MACRO RA1SHD512X64
  PIN A[0]
    AntennaGateArea  0.0792 ;
  END A[0]
  PIN A[1]
    AntennaGateArea  0.0792 ;
  END A[1]
  PIN A[2]
    AntennaGateArea  0.0792 ;
  END A[2]
  PIN A[3]
    AntennaGateArea  0.0792 ;
  END A[3]
  PIN A[4]
    AntennaGateArea  0.0792 ;
  END A[4]
  PIN A[5]
    AntennaGateArea  0.0792 ;
  END A[5]
  PIN A[6]
    AntennaGateArea  0.0792 ;
  END A[6]
  PIN A[7]
    AntennaGateArea  0.0792 ;
  END A[7]
  PIN A[8]
    AntennaGateArea  0.0792 ;
  END A[8]
  PIN CEN
    AntennaGateArea  0.0792 ;
  END CEN
  PIN CLK
    AntennaGateArea  0.0792 ;
  END CLK
  PIN D[0]
    AntennaGateArea  0.0792 ;
  END D[0]
  PIN D[10]
    AntennaGateArea  0.0792 ;
  END D[10]
  PIN D[11]
    AntennaGateArea  0.0792 ;
  END D[11]
  PIN D[12]
    AntennaGateArea  0.0792 ;
  END D[12]
  PIN D[13]
    AntennaGateArea  0.0792 ;
  END D[13]
  PIN D[14]
    AntennaGateArea  0.0792 ;
  END D[14]
  PIN D[15]
    AntennaGateArea  0.0792 ;
  END D[15]
  PIN D[16]
    AntennaGateArea  0.0792 ;
  END D[16]
  PIN D[17]
    AntennaGateArea  0.0792 ;
  END D[17]
  PIN D[18]
    AntennaGateArea  0.0792 ;
  END D[18]
  PIN D[19]
    AntennaGateArea  0.0792 ;
  END D[19]
  PIN D[1]
    AntennaGateArea  0.0792 ;
  END D[1]
  PIN D[20]
    AntennaGateArea  0.0792 ;
  END D[20]
  PIN D[21]
    AntennaGateArea  0.0792 ;
  END D[21]
  PIN D[22]
    AntennaGateArea  0.0792 ;
  END D[22]
  PIN D[23]
    AntennaGateArea  0.0792 ;
  END D[23]
  PIN D[24]
    AntennaGateArea  0.0792 ;
  END D[24]
  PIN D[25]
    AntennaGateArea  0.0792 ;
  END D[25]
  PIN D[26]
    AntennaGateArea  0.0792 ;
  END D[26]
  PIN D[27]
    AntennaGateArea  0.0792 ;
  END D[27]
  PIN D[28]
    AntennaGateArea  0.0792 ;
  END D[28]
  PIN D[29]
    AntennaGateArea  0.0792 ;
  END D[29]
  PIN D[2]
    AntennaGateArea  0.0792 ;
  END D[2]
  PIN D[30]
    AntennaGateArea  0.0792 ;
  END D[30]
  PIN D[31]
    AntennaGateArea  0.0792 ;
  END D[31]
  PIN D[32]
    AntennaGateArea  0.0792 ;
  END D[32]
  PIN D[33]
    AntennaGateArea  0.0792 ;
  END D[33]
  PIN D[34]
    AntennaGateArea  0.0792 ;
  END D[34]
  PIN D[35]
    AntennaGateArea  0.0792 ;
  END D[35]
  PIN D[36]
    AntennaGateArea  0.0792 ;
  END D[36]
  PIN D[37]
    AntennaGateArea  0.0792 ;
  END D[37]
  PIN D[38]
    AntennaGateArea  0.0792 ;
  END D[38]
  PIN D[39]
    AntennaGateArea  0.0792 ;
  END D[39]
  PIN D[3]
    AntennaGateArea  0.0792 ;
  END D[3]
  PIN D[40]
    AntennaGateArea  0.0792 ;
  END D[40]
  PIN D[41]
    AntennaGateArea  0.0792 ;
  END D[41]
  PIN D[42]
    AntennaGateArea  0.0792 ;
  END D[42]
  PIN D[43]
    AntennaGateArea  0.0792 ;
  END D[43]
  PIN D[44]
    AntennaGateArea  0.0792 ;
  END D[44]
  PIN D[45]
    AntennaGateArea  0.0792 ;
  END D[45]
  PIN D[46]
    AntennaGateArea  0.0792 ;
  END D[46]
  PIN D[47]
    AntennaGateArea  0.0792 ;
  END D[47]
  PIN D[48]
    AntennaGateArea  0.0792 ;
  END D[48]
  PIN D[49]
    AntennaGateArea  0.0792 ;
  END D[49]
  PIN D[4]
    AntennaGateArea  0.0792 ;
  END D[4]
  PIN D[50]
    AntennaGateArea  0.0792 ;
  END D[50]
  PIN D[51]
    AntennaGateArea  0.0792 ;
  END D[51]
  PIN D[52]
    AntennaGateArea  0.0792 ;
  END D[52]
  PIN D[53]
    AntennaGateArea  0.0792 ;
  END D[53]
  PIN D[54]
    AntennaGateArea  0.0792 ;
  END D[54]
  PIN D[55]
    AntennaGateArea  0.0792 ;
  END D[55]
  PIN D[56]
    AntennaGateArea  0.0792 ;
  END D[56]
  PIN D[57]
    AntennaGateArea  0.0792 ;
  END D[57]
  PIN D[58]
    AntennaGateArea  0.0792 ;
  END D[58]
  PIN D[59]
    AntennaGateArea  0.0792 ;
  END D[59]
  PIN D[5]
    AntennaGateArea  0.0792 ;
  END D[5]
  PIN D[60]
    AntennaGateArea  0.0792 ;
  END D[60]
  PIN D[61]
    AntennaGateArea  0.0792 ;
  END D[61]
  PIN D[62]
    AntennaGateArea  0.0792 ;
  END D[62]
  PIN D[63]
    AntennaGateArea  0.0792 ;
  END D[63]
  PIN D[6]
    AntennaGateArea  0.0792 ;
  END D[6]
  PIN D[7]
    AntennaGateArea  0.0792 ;
  END D[7]
  PIN D[8]
    AntennaGateArea  0.0792 ;
  END D[8]
  PIN D[9]
    AntennaGateArea  0.0792 ;
  END D[9]
  PIN OEN
    AntennaGateArea  0.0792 ;
  END OEN
  PIN WEN[0]
    AntennaGateArea  0.0792 ;
  END WEN[0]
  PIN WEN[1]
    AntennaGateArea  0.0792 ;
  END WEN[1]
  PIN WEN[2]
    AntennaGateArea  0.0792 ;
  END WEN[2]
  PIN WEN[3]
    AntennaGateArea  0.0792 ;
  END WEN[3]
  PIN WEN[4]
    AntennaGateArea  0.0792 ;
  END WEN[4]
  PIN WEN[5]
    AntennaGateArea  0.0792 ;
  END WEN[5]
  PIN WEN[6]
    AntennaGateArea  0.0792 ;
  END WEN[6]
  PIN WEN[7]
    AntennaGateArea  0.0792 ;
  END WEN[7]
END RA1SHD512X64
