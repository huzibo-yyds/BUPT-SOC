.SUBCKT AD1UHDV1 A B CI CO S VDD VSS VNW VPW
MM27 CO net111 VDD VNW p18 W=0.95u L=180.00n
MM25 S net79 VDD VNW p18 W=1.01u L=180.00n
MM23 net31 CI VDD VNW p18 W=580.0n L=180.00n
MM19 net31 A VDD VNW p18 W=0.545u L=180.00n
MM18 net31 B VDD VNW p18 W=580.0n L=180.00n
MM17 net79 net111 net31 VNW p18 W=580.0n L=180.00n
MM15 net18 CI VDD VNW p18 W=580.0n L=180.00n
MM12 net22 B net18 VNW p18 W=580.0n L=180.00n
MM11 net79 A net22 VNW p18 W=0.44u L=180.00n
MM8 net111 A net42 VNW p18 W=0.49u L=180.00n
MM7 net42 B VDD VNW p18 W=580.0n L=180.00n
MM4 net111 CI net55 VNW p18 W=580.0n L=180.00n
MM3 net55 B VDD VNW p18 W=580.0n L=180.00n
MM1 net55 A VDD VNW p18 W=580.0n L=180.00n
MM28 CO net111 VSS VPW n18 W=720.00n L=180.00n
MM26 S net79 VSS VPW n18 W=720.00n L=180.00n
MM24 net91 CI VSS VPW n18 W=430.00n L=180.00n
MM22 net79 net111 net91 VPW n18 W=430.00n L=180.00n
MM21 net91 B VSS VPW n18 W=430.00n L=180.00n
MM20 net91 A VSS VPW n18 W=430.00n L=180.00n
MM16 net67 CI VSS VPW n18 W=430.00n L=180.00n
MM14 net71 B net67 VPW n18 W=340.00n L=180.00n
MM13 net79 A net71 VPW n18 W=340.00n L=180.00n
MM10 net111 A net99 VPW n18 W=340.00n L=180.00n
MM9 net99 B VSS VPW n18 W=340.00n L=180.00n
MM6 net111 CI net103 VPW n18 W=430.00n L=180.00n
MM5 net103 B VSS VPW n18 W=430.00n L=180.00n
MM2 net103 A VSS VPW n18 W=0.42u L=180.00n
.ENDS AD1UHDV1
.SUBCKT AD1UHDV2 A B CI CO S VDD VSS VNW VPW
MM6 net3 CI net11 VPW n18 W=630.00n L=180.00n
MM5 net11 B VSS VPW n18 W=0.5u L=180.00n
MM2 net11 A VSS VPW n18 W=720.00n L=180.00n
MM9 net15 B VSS VPW n18 W=0.5u L=180.00n
MM10 net3 A net15 VPW n18 W=800.00n L=180.00n
MM20 net23 A VSS VPW n18 W=720.00n L=180.00n
MM21 net23 B VSS VPW n18 W=720.00n L=180.00n
MM24 net23 CI VSS VPW n18 W=540.00n L=180.00n
MM22 net35 net3 net23 VPW n18 W=720.00n L=180.00n
MM13 net35 A net43 VPW n18 W=400.00n L=180.00n
MM14 net43 B net47 VPW n18 W=400.00n L=180.00n
MM16 net47 CI VSS VPW n18 W=770.00n L=180.00n
MM26 S net35 VSS VPW n18 W=1.44u L=180.00n
MM28 CO net3 VSS VPW n18 W=1.44u L=180.00n
MM1 net59 A VDD VNW p18 W=990.0n L=180.00n
MM3 net59 B VDD VNW p18 W=0.69u L=180.00n
MM4 net3 CI net59 VNW p18 W=990.0n L=180.00n
MM7 net78 B VDD VNW p18 W=720.0n L=180.00n
MM8 net3 A net78 VNW p18 W=490.0n L=180.00n
MM18 net83 B VDD VNW p18 W=0.58u L=180.00n
MM19 net83 A VDD VNW p18 W=0.545u L=180.00n
MM23 net83 CI VDD VNW p18 W=0.98u L=180.00n
MM17 net35 net3 net83 VNW p18 W=0.95u L=180.00n
MM11 net35 A net98 VNW p18 W=0.44u L=180.00n
MM12 net98 B net102 VNW p18 W=0.83u L=180.00n
MM15 net102 CI VDD VNW p18 W=0.85u L=180.00n
MM25 S net35 VDD VNW p18 W=2.02u L=180.00n
MM27 CO net3 VDD VNW p18 W=2.02u L=180.00n
.ENDS AD1UHDV2
.SUBCKT ADH1UHDV1 A B CO S VDD VSS VNW VPW
MM12 S net053 VSS VPW n18 W=720.00n L=180.00n
MM11 net056 net20 VSS VPW n18 W=0.72u L=180.00n
MM5 net053 B net056 VPW n18 W=0.385u L=180.00n
MM4 net053 A net056 VPW n18 W=0.385u L=180.00n
MM2 CO net20 VSS VPW n18 W=720.00n L=180.00n
MM9 net8 B VSS VPW n18 W=0.475u L=180.00n
MM10 net20 A net8 VPW n18 W=0.475u L=180.00n
MM6 net053 net20 VDD VNW p18 W=0.595u L=180.00n
MM7 net080 A VDD VNW p18 W=0.595u L=180.00n
MM13 S net053 VDD VNW p18 W=1.01u L=180.00n
MM8 net053 B net080 VNW p18 W=0.595u L=180.00n
MM0 CO net20 VDD VNW p18 W=1.01u L=180.00n
MM1 net20 A VDD VNW p18 W=0.595u L=180.00n
MM3 net20 B VDD VNW p18 W=0.595u L=180.00n
.ENDS ADH1UHDV1
.SUBCKT ADH1UHDV2 A B CO S VDD VSS VNW VPW
MM3 net9 B VDD VNW p18 W=0.97u L=180.00n
MM1 net9 A VDD VNW p18 W=0.97u L=180.00n
MM0 CO net9 VDD VNW p18 W=2.02u L=180.00n
MM6 net45 net9 VDD VNW p18 W=0.65u L=180.00n
MM8 net45 B net24 VNW p18 W=950.0n L=180.00n
MM7 net24 A VDD VNW p18 W=950.0n L=180.00n
MM13 S net45 VDD VNW p18 W=2.02u L=180.00n
MM10 net9 A net37 VPW n18 W=0.635u L=180.00n
MM9 net37 B VSS VPW n18 W=0.635u L=180.00n
MM2 CO net9 VSS VPW n18 W=1.36u L=180.00n
MM4 net45 A net48 VPW n18 W=0.635u L=180.00n
MM5 net45 B net48 VPW n18 W=0.635u L=180.00n
MM11 net48 net9 VSS VPW n18 W=0.635u L=180.00n
MM12 S net45 VSS VPW n18 W=1.44u L=180.00n
.ENDS ADH1UHDV2
.SUBCKT ADH1UHDV3 A B CO S VDD VSS VNW VPW
MM12 S net17 VSS VPW n18 W=2.16u L=180.00n
MM11 net20 net53 VSS VPW n18 W=720.00n L=180.00n
MM5 net17 B net20 VPW n18 W=720.00n L=180.00n
MM4 net17 A net20 VPW n18 W=720.00n L=180.00n
MM2 CO net53 VSS VPW n18 W=2.16u L=180.00n
MM9 net25 B VSS VPW n18 W=720.00n L=180.00n
MM10 net53 A net25 VPW n18 W=720.00n L=180.00n
MM13 S net17 VDD VNW p18 W=3.03u L=180.00n
MM7 net44 A VDD VNW p18 W=0.95u L=180.00n
MM8 net17 B net44 VNW p18 W=0.95u L=180.00n
MM6 net17 net53 VDD VNW p18 W=0.95u L=180.00n
MM0 CO net53 VDD VNW p18 W=3.03u L=180.00n
MM1 net53 A VDD VNW p18 W=0.97u L=180.00n
MM3 net53 B VDD VNW p18 W=0.97u L=180.00n
.ENDS ADH1UHDV3
.SUBCKT AND2UHDV0P4 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=0.28u L=180.00n
MM3 net24 A1 net8 VPW n18 W=0.28u L=180.00n
MM5 net8 A2 VSS VPW n18 W=0.28u L=180.00n
MM1 Z net24 VDD VNW p18 W=0.475u L=180.00n
MM0 net24 A2 VDD VNW p18 W=0.475u L=180.00n
MM2 net24 A1 VDD VNW p18 W=0.475u L=180.00n
.ENDS AND2UHDV0P4
****Sub-Circuit for AND2UHDV0P7, Tue Jun 13 18:01:17 CST 2017****
.SUBCKT AND2UHDV0P7 A1 A2 Z VDD VSS VNW VPW
MM3 net4 A1 net20 VPW n18 W=475.00n L=180.00n
MM5 net20 A2 VSS VPW n18 W=475.00n L=180.00n
MM4 Z net4 VSS VPW n18 W=560.00n L=180.00n
MM2 net4 A1 VDD VNW p18 W=475.00n L=180.00n
MM0 net4 A2 VDD VNW p18 W=475.00n L=180.00n
MM1 Z net4 VDD VNW p18 W=790.00n L=180.00n
.ENDS AND2UHDV0P7
.SUBCKT AND2UHDV1 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=720.00n L=180.00n
MM5 net8 A2 VSS VPW n18 W=0.475u L=180.00n
MM3 net24 A1 net8 VPW n18 W=0.475u L=180.00n
MM1 Z net24 VDD VNW p18 W=1.01u L=180.00n
MM0 net24 A2 VDD VNW p18 W=0.475u L=180.00n
MM2 net24 A1 VDD VNW p18 W=0.515u L=180.00n
.ENDS AND2UHDV1
.SUBCKT AND2UHDV2 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=1.44u L=180.00n
MM5 net8 A2 VSS VPW n18 W=720.00n L=180.00n
MM3 net24 A1 net8 VPW n18 W=720.00n L=180.00n
MM1 Z net24 VDD VNW p18 W=2.02u L=180.00n
MM0 net24 A2 VDD VNW p18 W=0.97u L=180.00n
MM2 net24 A1 VDD VNW p18 W=0.97u L=180.00n
.ENDS AND2UHDV2
.SUBCKT AND2UHDV3 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=2.16u L=180.00n
MM5 net8 A2 VSS VPW n18 W=720.00n L=180.00n
MM3 net24 A1 net8 VPW n18 W=720.00n L=180.00n
MM1 Z net24 VDD VNW p18 W=3.03u L=180.00n
MM0 net24 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net24 A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS AND2UHDV3
.SUBCKT AND2UHDV4 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=2.88u L=180.00n
MM5 net8 A2 VSS VPW n18 W=1.15u L=180.00n
MM3 net24 A1 net8 VPW n18 W=1.15u L=180.00n
MM1 Z net24 VDD VNW p18 W=4.04u L=180.00n
MM0 net24 A2 VDD VNW p18 W=1.52u L=180.00n
MM2 net24 A1 VDD VNW p18 W=1.52u L=180.00n
.ENDS AND2UHDV4
.SUBCKT AND2UHDV6 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=4.32u L=180.00n
MM5 net8 A2 VSS VPW n18 W=1.44u L=180.00n
MM3 net24 A1 net8 VPW n18 W=1.44u L=180.00n
MM1 Z net24 VDD VNW p18 W=6.06u L=180.00n
MM0 net24 A2 VDD VNW p18 W=2.02u L=180.00n
MM2 net24 A1 VDD VNW p18 W=2.02u L=180.00n
.ENDS AND2UHDV6
.SUBCKT AND2UHDV8 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=5.76u L=180.00n
MM5 net8 A2 VSS VPW n18 W=2.16u L=180.00n
MM3 net24 A1 net8 VPW n18 W=2.16u L=180.00n
MM1 Z net24 VDD VNW p18 W=8.08u L=180.00n
MM0 net24 A2 VDD VNW p18 W=3.03u L=180.00n
MM2 net24 A1 VDD VNW p18 W=3.03u L=180.00n
.ENDS AND2UHDV8
.SUBCKT AND3UHDV0P7 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net5 A3 VSS VPW n18 W=0.475u L=180.00n
MM4 Z net33 VSS VPW n18 W=0.605u L=180.00n
MM5 net13 A2 net5 VPW n18 W=0.475u L=180.00n
MM3 net33 A1 net13 VPW n18 W=0.475u L=180.00n
MM6 net33 A3 VDD VNW p18 W=0.51u L=180.00n
MM1 Z net33 VDD VNW p18 W=0.8u L=180.00n
MM0 net33 A2 VDD VNW p18 W=0.51u L=180.00n
MM2 net33 A1 VDD VNW p18 W=0.51u L=180.00n
.ENDS AND3UHDV0P7
.SUBCKT AND3UHDV1 A1 A2 A3 Z VDD VSS VNW VPW
MM2 net5 A1 VDD VNW p18 W=0.575u L=180.00n
MM0 net5 A2 VDD VNW p18 W=0.575u L=180.00n
MM1 Z net5 VDD VNW p18 W=1.01u L=180.00n
MM6 net5 A3 VDD VNW p18 W=0.575u L=180.00n
MM3 net5 A1 net25 VPW n18 W=0.475u L=180.00n
MM5 net25 A2 net33 VPW n18 W=0.475u L=180.00n
MM4 Z net5 VSS VPW n18 W=720.00n L=180.00n
MM7 net33 A3 VSS VPW n18 W=0.475u L=180.00n
.ENDS AND3UHDV1
.SUBCKT AND3UHDV2 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net5 A3 VSS VPW n18 W=720.00n L=180.00n
MM4 Z net33 VSS VPW n18 W=1.44u L=180.00n
MM5 net13 A2 net5 VPW n18 W=720.00n L=180.00n
MM3 net33 A1 net13 VPW n18 W=720.00n L=180.00n
MM6 net33 A3 VDD VNW p18 W=0.97u L=180.00n
MM1 Z net33 VDD VNW p18 W=2.02u L=180.00n
MM0 net33 A2 VDD VNW p18 W=0.97u L=180.00n
MM2 net33 A1 VDD VNW p18 W=0.97u L=180.00n
.ENDS AND3UHDV2
.SUBCKT AND3UHDV3 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net5 A3 VSS VPW n18 W=720.00n L=180.00n
MM4 Z net33 VSS VPW n18 W=2.16u L=180.00n
MM5 net13 A2 net5 VPW n18 W=720.00n L=180.00n
MM3 net33 A1 net13 VPW n18 W=720.00n L=180.00n
MM6 net33 A3 VDD VNW p18 W=1.01u L=180.00n
MM1 Z net33 VDD VNW p18 W=3.03u L=180.00n
MM0 net33 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net33 A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS AND3UHDV3
.SUBCKT AND3UHDV4 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net5 A3 VSS VPW n18 W=1.01u L=180.00n
MM4 Z net33 VSS VPW n18 W=2.88u L=180.00n
MM5 net13 A2 net5 VPW n18 W=1.01u L=180.00n
MM3 net33 A1 net13 VPW n18 W=1.01u L=180.00n
MM6 net33 A3 VDD VNW p18 W=1.51u L=180.00n
MM1 Z net33 VDD VNW p18 W=4.04u L=180.00n
MM0 net33 A2 VDD VNW p18 W=1.51u L=180.00n
MM2 net33 A1 VDD VNW p18 W=1.51u L=180.00n
.ENDS AND3UHDV4
.SUBCKT AND4UHDV0P7 A1 A2 A3 A4 Z VDD VSS VNW VPW
MM8 net14 A4 VDD VNW p18 W=0.51u L=180.00n
MM2 net14 A1 VDD VNW p18 W=0.51u L=180.00n
MM0 net14 A2 VDD VNW p18 W=0.51u L=180.00n
MM1 Z net14 VDD VNW p18 W=0.8u L=180.00n
MM6 net14 A3 VDD VNW p18 W=0.51u L=180.00n
MM9 net30 A4 VSS VPW n18 W=0.475u L=180.00n
MM3 net14 A1 net38 VPW n18 W=0.475u L=180.00n
MM5 net38 A2 net42 VPW n18 W=0.475u L=180.00n
MM4 Z net14 VSS VPW n18 W=0.605u L=180.00n
MM7 net42 A3 net30 VPW n18 W=0.475u L=180.00n
.ENDS AND4UHDV0P7
.SUBCKT AND4UHDV1 A1 A2 A3 A4 Z VDD VSS VNW VPW
MM7 net6 A3 net18 VPW n18 W=0.475u L=180.00n
MM5 net10 A2 net6 VPW n18 W=0.475u L=180.00n
MM3 net34 A1 net10 VPW n18 W=0.475u L=180.00n
MM9 net18 A4 VSS VPW n18 W=0.475u L=180.00n
MM4 Z net34 VSS VPW n18 W=720.00n L=180.00n
MM6 net34 A3 VDD VNW p18 W=0.575u L=180.00n
MM0 net34 A2 VDD VNW p18 W=0.575u L=180.00n
MM2 net34 A1 VDD VNW p18 W=0.575u L=180.00n
MM8 net34 A4 VDD VNW p18 W=0.575u L=180.00n
MM1 Z net34 VDD VNW p18 W=1.01u L=180.00n
.ENDS AND4UHDV1
.SUBCKT AND4UHDV2 A1 A2 A3 A4 Z VDD VSS VNW VPW
MM7 net6 A3 net18 VPW n18 W=0.675u L=180.00n
MM5 net10 A2 net6 VPW n18 W=0.675u L=180.00n
MM3 net34 A1 net10 VPW n18 W=0.675u L=180.00n
MM9 net18 A4 VSS VPW n18 W=0.675u L=180.00n
MM4 Z net34 VSS VPW n18 W=1.44u L=180.00n
MM6 net34 A3 VDD VNW p18 W=0.89u L=180.00n
MM0 net34 A2 VDD VNW p18 W=0.89u L=180.00n
MM2 net34 A1 VDD VNW p18 W=0.89u L=180.00n
MM8 net34 A4 VDD VNW p18 W=0.89u L=180.00n
MM1 Z net34 VDD VNW p18 W=2.02u L=180.00n
.ENDS AND4UHDV2
.SUBCKT AND4UHDV3 A1 A2 A3 A4 Z VDD VSS VNW VPW
MM7 net6 A3 net18 VPW n18 W=0.675u L=180.00n
MM5 net10 A2 net6 VPW n18 W=0.675u L=180.00n
MM3 net34 A1 net10 VPW n18 W=0.675u L=180.00n
MM9 net18 A4 VSS VPW n18 W=0.675u L=180.00n
MM4 Z net34 VSS VPW n18 W=2.16u L=180.00n
MM6 net34 A3 VDD VNW p18 W=0.89u L=180.00n
MM0 net34 A2 VDD VNW p18 W=0.89u L=180.00n
MM2 net34 A1 VDD VNW p18 W=0.89u L=180.00n
MM8 net34 A4 VDD VNW p18 W=0.89u L=180.00n
MM1 Z net34 VDD VNW p18 W=3.03u L=180.00n
.ENDS AND4UHDV3
.SUBCKT AO112UHDV0P4 A1 A2 B C Z VDD VSS VNW VPW
MM7 net17 B VDD VNW p18 W=0.495u L=180.00n
MM6 net21 C net17 VNW p18 W=0.495u L=180.00n
MM2 net18 A1 net21 VNW p18 W=0.495u L=180.00n
MM0 net18 A2 net21 VNW p18 W=0.495u L=180.00n
MM1 Z net18 VDD VNW p18 W=0.495u L=180.00n
MM9 net18 B VSS VPW n18 W=0.275u L=180.00n
MM8 net18 C VSS VPW n18 W=0.275u L=180.00n
MM5 net38 A2 VSS VPW n18 W=0.28u L=180.00n
MM3 net18 A1 net38 VPW n18 W=0.28u L=180.00n
MM4 Z net18 VSS VPW n18 W=0.28u L=180.00n
.ENDS AO112UHDV0P4
.SUBCKT AO112UHDV0P7 A1 A2 B C Z VDD VSS VNW VPW
MM3 net30 A1 net10 VPW n18 W=0.42u L=180.00n
MM5 net10 A2 VSS VPW n18 W=0.42u L=180.00n
MM8 net30 C VSS VPW n18 W=0.42u L=180.00n
MM9 net30 B VSS VPW n18 W=0.42u L=180.00n
MM4 Z net30 VSS VPW n18 W=560.00n L=180.00n
MM0 net30 A2 net33 VNW p18 W=0.495u L=180.00n
MM2 net30 A1 net33 VNW p18 W=0.495u L=180.00n
MM6 net33 C net37 VNW p18 W=0.495u L=180.00n
MM7 net37 B VDD VNW p18 W=0.495u L=180.00n
MM1 Z net30 VDD VNW p18 W=790.0n L=180.00n
.ENDS AO112UHDV0P7
.SUBCKT AO112UHDV1 A1 A2 B C Z VDD VSS VNW VPW
MM3 net30 A1 net10 VPW n18 W=0.42u L=180.00n
MM5 net10 A2 VSS VPW n18 W=0.42u L=180.00n
MM8 net30 C VSS VPW n18 W=0.42u L=180.00n
MM9 net30 B VSS VPW n18 W=0.42u L=180.00n
MM4 Z net30 VSS VPW n18 W=0.695u L=180.00n
MM0 net30 A2 net33 VNW p18 W=0.495u L=180.00n
MM2 net30 A1 net33 VNW p18 W=0.495u L=180.00n
MM6 net33 C net37 VNW p18 W=0.56u L=180.00n
MM7 net37 B VDD VNW p18 W=0.56u L=180.00n
MM1 Z net30 VDD VNW p18 W=0.915u L=180.00n
.ENDS AO112UHDV1
.SUBCKT AO112UHDV2 A1 A2 B C Z VDD VSS VNW VPW
MM3 net30 A1 net10 VPW n18 W=0.62u L=180.00n
MM5 net10 A2 VSS VPW n18 W=0.62u L=180.00n
MM8 net30 C VSS VPW n18 W=0.62u L=180.00n
MM9 net30 B VSS VPW n18 W=0.62u L=180.00n
MM4 Z net30 VSS VPW n18 W=1.44u L=180.00n
MM0 net30 A2 net33 VNW p18 W=0.97u L=180.00n
MM2 net30 A1 net33 VNW p18 W=0.97u L=180.00n
MM6 net33 C net37 VNW p18 W=0.97u L=180.00n
MM7 net37 B VDD VNW p18 W=0.97u L=180.00n
MM1 Z net30 VDD VNW p18 W=2.02u L=180.00n
.ENDS AO112UHDV2
.SUBCKT AO112UHDV3 A1 A2 B C Z VDD VSS VNW VPW
MM3 net30 A1 net10 VPW n18 W=720.00n L=180.00n
MM5 net10 A2 VSS VPW n18 W=720.00n L=180.00n
MM8 net30 C VSS VPW n18 W=720.00n L=180.00n
MM9 net30 B VSS VPW n18 W=720.00n L=180.00n
MM4 Z net30 VSS VPW n18 W=2.16u L=180.00n
MM0 net30 A2 net33 VNW p18 W=1.01u L=180.00n
MM2 net30 A1 net33 VNW p18 W=1.01u L=180.00n
MM6 net33 C net37 VNW p18 W=1.01u L=180.00n
MM7 net37 B VDD VNW p18 W=1.01u L=180.00n
MM1 Z net30 VDD VNW p18 W=3.03u L=180.00n
.ENDS AO112UHDV3
.SUBCKT AO12UHDV0P4 A1 A2 B Z VDD VSS VNW VPW
MM4 Z net33 VSS VPW n18 W=430.00n L=180.00n
MM3 net33 A1 net13 VPW n18 W=430.00n L=180.00n
MM5 net13 A2 VSS VPW n18 W=430.00n L=180.00n
MM8 net33 B VSS VPW n18 W=430.00n L=180.00n
MM1 Z net33 VDD VNW p18 W=490.0n L=180.00n
MM0 net33 A2 net36 VNW p18 W=490.0n L=180.00n
MM2 net33 A1 net36 VNW p18 W=490.0n L=180.00n
MM7 net36 B VDD VNW p18 W=490.0n L=180.00n
.ENDS AO12UHDV0P4
.SUBCKT AO12UHDV0P7 A1 A2 B Z VDD VSS VNW VPW
MM2 net5 A1 net8 VNW p18 W=500.0n L=180.00n
MM0 net5 A2 net8 VNW p18 W=500.0n L=180.00n
MM7 net8 B VDD VNW p18 W=500.0n L=180.00n
MM1 Z net5 VDD VNW p18 W=790.0n L=180.00n
MM8 net5 B VSS VPW n18 W=430.00n L=180.00n
MM5 net25 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 net5 A1 net25 VPW n18 W=430.00n L=180.00n
MM4 Z net5 VSS VPW n18 W=560.00n L=180.00n
.ENDS AO12UHDV0P7
.SUBCKT AO12UHDV1 A1 A2 B Z VDD VSS VNW VPW
MM2 net5 A1 net8 VNW p18 W=580.0n L=180.00n
MM0 net5 A2 net8 VNW p18 W=580.0n L=180.00n
MM7 net8 B VDD VNW p18 W=580.0n L=180.00n
MM1 Z net5 VDD VNW p18 W=0.92u L=180.00n
MM8 net5 B VSS VPW n18 W=430.00n L=180.00n
MM5 net25 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 net5 A1 net25 VPW n18 W=430.00n L=180.00n
MM4 Z net5 VSS VPW n18 W=720.00n L=180.00n
.ENDS AO12UHDV1
.SUBCKT AO12UHDV2 A1 A2 B Z VDD VSS VNW VPW
MM2 net5 A1 net8 VNW p18 W=950.0n L=180.00n
MM0 net5 A2 net8 VNW p18 W=950.0n L=180.00n
MM7 net8 B VDD VNW p18 W=950.0n L=180.00n
MM1 Z net5 VDD VNW p18 W=2.02u L=180.00n
MM8 net5 B VSS VPW n18 W=630.00n L=180.00n
MM5 net25 A2 VSS VPW n18 W=630.00n L=180.00n
MM3 net5 A1 net25 VPW n18 W=630.00n L=180.00n
MM4 Z net5 VSS VPW n18 W=1.44u L=180.00n
.ENDS AO12UHDV2
.SUBCKT AO12UHDV3 A1 A2 B Z VDD VSS VNW VPW
MM2 net5 A1 net8 VNW p18 W=1.01u L=180.00n
MM0 net5 A2 net8 VNW p18 W=1.01u L=180.00n
MM7 net8 B VDD VNW p18 W=1.01u L=180.00n
MM1 Z net5 VDD VNW p18 W=3.03u L=180.00n
MM8 net5 B VSS VPW n18 W=720.00n L=180.00n
MM5 net25 A2 VSS VPW n18 W=720.00n L=180.00n
MM3 net5 A1 net25 VPW n18 W=720.00n L=180.00n
MM4 Z net5 VSS VPW n18 W=2.16u L=180.00n
.ENDS AO12UHDV3
.SUBCKT AO12UHDV4 A1 A2 B Z VDD VSS VNW VPW
MM2 net5 A1 net8 VNW p18 W=1.35u L=180.00n
MM0 net5 A2 net8 VNW p18 W=1.35u L=180.00n
MM7 net8 B VDD VNW p18 W=1.35u L=180.00n
MM1 Z net5 VDD VNW p18 W=4.04u L=180.00n
MM8 net5 B VSS VPW n18 W=1060.00n L=180.00n
MM5 net25 A2 VSS VPW n18 W=1060.00n L=180.00n
MM3 net5 A1 net25 VPW n18 W=1060.00n L=180.00n
MM4 Z net5 VSS VPW n18 W=2.88u L=180.00n
.ENDS AO12UHDV4
.SUBCKT AO21BUHDV0P4 A1 A2 B Z VDD VSS VNW VPW
MM3 Z B net9 VPW n18 W=0.28u L=180.00n
MM1 net9 net044 VSS VPW n18 W=0.28u L=180.00n
MM6 net13 A2 VSS VPW n18 W=0.28u L=180.00n
MM9 net044 A1 net13 VPW n18 W=0.28u L=180.00n
MM5 Z net044 VDD VNW p18 W=0.425u L=180.00n
MM4 Z B VDD VNW p18 W=0.425u L=180.00n
MM0 net044 A1 VDD VNW p18 W=0.425u L=180.00n
MM2 net044 A2 VDD VNW p18 W=0.425u L=180.00n
.ENDS AO21BUHDV0P4
.SUBCKT AO21BUHDV0P7 A1 A2 B Z VDD VSS VNW VPW
MM5 Z net16 VDD VNW p18 W=790.0n L=180.00n
MM4 Z B VDD VNW p18 W=790.0n L=180.00n
MM0 net16 A1 VDD VNW p18 W=500.0n L=180.00n
MM2 net16 A2 VDD VNW p18 W=500.0n L=180.00n
MM3 Z B net40 VPW n18 W=560.00n L=180.00n
MM1 net40 net16 VSS VPW n18 W=560.00n L=180.00n
MM6 net36 A2 VSS VPW n18 W=430.00n L=180.00n
MM9 net16 A1 net36 VPW n18 W=430.00n L=180.00n
.ENDS AO21BUHDV0P7
.SUBCKT AO21BUHDV1 A1 A2 B Z VDD VSS VNW VPW
MM5 Z net16 VDD VNW p18 W=1.01u L=180.00n
MM4 Z B VDD VNW p18 W=1.01u L=180.00n
MM0 net16 A1 VDD VNW p18 W=580.0n L=180.00n
MM2 net16 A2 VDD VNW p18 W=580.0n L=180.00n
MM3 Z B net40 VPW n18 W=720.00n L=180.00n
MM1 net40 net16 VSS VPW n18 W=720.00n L=180.00n
MM6 net36 A2 VSS VPW n18 W=430.00n L=180.00n
MM9 net16 A1 net36 VPW n18 W=430.00n L=180.00n
.ENDS AO21BUHDV1
.SUBCKT AO21BUHDV2 A1 A2 B Z VDD VSS VNW VPW
MM5 Z net16 VDD VNW p18 W=2.02u L=180.00n
MM4 Z B VDD VNW p18 W=1.9u L=180.00n
MM0 net16 A1 VDD VNW p18 W=950.0n L=180.00n
MM2 net16 A2 VDD VNW p18 W=950.0n L=180.00n
MM3 Z B net40 VPW n18 W=1.44u L=180.00n
MM1 net40 net16 VSS VPW n18 W=1.44u L=180.00n
MM6 net36 A2 VSS VPW n18 W=630.00n L=180.00n
MM9 net16 A1 net36 VPW n18 W=630.00n L=180.00n
.ENDS AO21BUHDV2
.SUBCKT AO21BUHDV3 A1 A2 B Z VDD VSS VNW VPW
MM5 Z net16 VDD VNW p18 W=2.97u L=180.00n
MM4 Z B VDD VNW p18 W=2.91u L=180.00n
MM0 net16 A1 VDD VNW p18 W=1.01u L=180.00n
MM2 net16 A2 VDD VNW p18 W=1.01u L=180.00n
MM3 Z B net40 VPW n18 W=2.16u L=180.00n
MM1 net40 net16 VSS VPW n18 W=2.16u L=180.00n
MM6 net36 A2 VSS VPW n18 W=720.00n L=180.00n
MM9 net16 A1 net36 VPW n18 W=720.00n L=180.00n
.ENDS AO21BUHDV3
.SUBCKT AO221UHDV0P4 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM11 net7 B2 VSS VPW n18 W=0.28u L=180.00n
MM3 net11 A1 net15 VPW n18 W=0.28u L=180.00n
MM5 net15 A2 VSS VPW n18 W=0.28u L=180.00n
MM8 net11 B1 net7 VPW n18 W=0.28u L=180.00n
MM9 net11 C VSS VPW n18 W=0.28u L=180.00n
MM4 Z net11 VSS VPW n18 W=0.28u L=180.00n
MM10 net35 B1 net38 VNW p18 W=0.495u L=180.00n
MM0 net38 A2 VDD VNW p18 W=0.5u L=180.00n
MM2 net38 A1 VDD VNW p18 W=0.5u L=180.00n
MM7 net11 C net35 VNW p18 W=0.485u L=180.00n
MM1 Z net11 VDD VNW p18 W=0.5u L=180.00n
MM6 net35 B2 net38 VNW p18 W=0.495u L=180.00n
.ENDS AO221UHDV0P4
.SUBCKT AO221UHDV0P7 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM1 Z net47 VDD VNW p18 W=790.0n L=180.00n
MM2 net26 A1 VDD VNW p18 W=500.0n L=180.00n
MM0 net26 A2 VDD VNW p18 W=500.0n L=180.00n
MM6 net23 B2 net26 VNW p18 W=0.495u L=180.00n
MM10 net23 B1 net26 VNW p18 W=0.495u L=180.00n
MM7 net47 C net23 VNW p18 W=0.485u L=180.00n
MM4 Z net47 VSS VPW n18 W=0.58u L=180.00n
MM9 net47 C VSS VPW n18 W=0.47u L=180.00n
MM8 net47 B1 net0134 VPW n18 W=0.47u L=180.00n
MM5 net43 A2 VSS VPW n18 W=0.47u L=180.00n
MM3 net47 A1 net43 VPW n18 W=0.47u L=180.00n
MM11 net0134 B2 VSS VPW n18 W=0.47u L=180.00n
.ENDS AO221UHDV0P7
.SUBCKT AO221UHDV1 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM1 Z net47 VDD VNW p18 W=1.01u L=180.00n
MM2 net26 A1 VDD VNW p18 W=580.0n L=180.00n
MM0 net26 A2 VDD VNW p18 W=580.0n L=180.00n
MM6 net23 B2 net26 VNW p18 W=580.0n L=180.00n
MM10 net23 B1 net26 VNW p18 W=580.0n L=180.00n
MM7 net47 C net23 VNW p18 W=580.0n L=180.00n
MM4 Z net47 VSS VPW n18 W=720.00n L=180.00n
MM9 net47 C VSS VPW n18 W=0.47u L=180.00n
MM8 net47 B1 net080 VPW n18 W=0.47u L=180.00n
MM5 net43 A2 VSS VPW n18 W=0.47u L=180.00n
MM3 net47 A1 net43 VPW n18 W=0.47u L=180.00n
MM11 net080 B2 VSS VPW n18 W=0.47u L=180.00n
.ENDS AO221UHDV1
.SUBCKT AO221UHDV2 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM1 Z net47 VDD VNW p18 W=2.02u L=180.00n
MM2 net26 A1 VDD VNW p18 W=0.97u L=180.00n
MM0 net26 A2 VDD VNW p18 W=0.97u L=180.00n
MM6 net23 B2 net26 VNW p18 W=0.97u L=180.00n
MM10 net23 B1 net26 VNW p18 W=0.97u L=180.00n
MM7 net47 C net23 VNW p18 W=0.97u L=180.00n
MM4 Z net47 VSS VPW n18 W=1.44u L=180.00n
MM9 net47 C VSS VPW n18 W=0.62u L=180.00n
MM8 net47 B1 net0134 VPW n18 W=0.62u L=180.00n
MM5 net43 A2 VSS VPW n18 W=0.62u L=180.00n
MM3 net47 A1 net43 VPW n18 W=0.62u L=180.00n
MM11 net0134 B2 VSS VPW n18 W=0.62u L=180.00n
.ENDS AO221UHDV2
.SUBCKT AO221UHDV3 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM1 Z net47 VDD VNW p18 W=3.03u L=180.00n
MM2 net26 A1 VDD VNW p18 W=1.01u L=180.00n
MM0 net26 A2 VDD VNW p18 W=1.01u L=180.00n
MM6 net23 B2 net26 VNW p18 W=1.01u L=180.00n
MM10 net23 B1 net26 VNW p18 W=1.01u L=180.00n
MM7 net47 C net23 VNW p18 W=1.01u L=180.00n
MM4 Z net47 VSS VPW n18 W=2.16u L=180.00n
MM9 net47 C VSS VPW n18 W=720.00n L=180.00n
MM8 net47 B1 net080 VPW n18 W=720.00n L=180.00n
MM5 net43 A2 VSS VPW n18 W=720.00n L=180.00n
MM3 net47 A1 net43 VPW n18 W=720.00n L=180.00n
MM11 net080 B2 VSS VPW n18 W=720.00n L=180.00n
.ENDS AO221UHDV3
.SUBCKT AO222UHDV0P4 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM16 net10 A1 net081 VPW n18 W=0.28u L=180.00n
MM15 net081 A2 VSS VPW n18 W=0.28u L=180.00n
MM4 Z net10 VSS VPW n18 W=0.28u L=180.00n
MM3 net10 B1 net14 VPW n18 W=0.28u L=180.00n
MM5 net14 B2 VSS VPW n18 W=0.28u L=180.00n
MM8 net10 C1 net085 VPW n18 W=0.28u L=180.00n
MM12 net085 C2 VSS VPW n18 W=0.28u L=180.00n
MM11 net0112 B1 net0116 VNW p18 W=490.0n L=180.00n
MM1 Z net10 VDD VNW p18 W=490.0n L=180.00n
MM6 net0116 A2 VDD VNW p18 W=490.0n L=180.00n
MM0 net10 C2 net0112 VNW p18 W=490.0n L=180.00n
MM2 net10 C1 net0112 VNW p18 W=490.0n L=180.00n
MM7 net0116 A1 VDD VNW p18 W=490.0n L=180.00n
MM10 net0112 B2 net0116 VNW p18 W=490.0n L=180.00n
.ENDS AO222UHDV0P4
.SUBCKT AO222UHDV0P7 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM1 Z net60 VDD VNW p18 W=790.0n L=180.00n
MM6 net27 A2 VDD VNW p18 W=500.0n L=180.00n
MM7 net27 A1 VDD VNW p18 W=500.0n L=180.00n
MM10 net31 B2 net27 VNW p18 W=500.0n L=180.00n
MM11 net31 B1 net27 VNW p18 W=500.0n L=180.00n
MM2 net60 C1 net31 VNW p18 W=500.0n L=180.00n
MM0 net60 C2 net31 VNW p18 W=500.0n L=180.00n
MM5 net36 B2 VSS VPW n18 W=430.00n L=180.00n
MM3 net60 B1 net36 VPW n18 W=430.00n L=180.00n
MM4 Z net60 VSS VPW n18 W=560.00n L=180.00n
MM8 net60 C1 net52 VPW n18 W=430.00n L=180.00n
MM12 net52 C2 VSS VPW n18 W=430.00n L=180.00n
MM15 net56 A2 VSS VPW n18 W=430.00n L=180.00n
MM16 net60 A1 net56 VPW n18 W=430.00n L=180.00n
.ENDS AO222UHDV0P7
.SUBCKT AO222UHDV1 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM1 Z net60 VDD VNW p18 W=0.98u L=180.00n
MM6 net27 A2 VDD VNW p18 W=580.0n L=180.00n
MM7 net27 A1 VDD VNW p18 W=580.0n L=180.00n
MM10 net31 B2 net27 VNW p18 W=580.0n L=180.00n
MM11 net31 B1 net27 VNW p18 W=580.0n L=180.00n
MM2 net60 C1 net31 VNW p18 W=580.0n L=180.00n
MM0 net60 C2 net31 VNW p18 W=580.0n L=180.00n
MM5 net36 B2 VSS VPW n18 W=430.00n L=180.00n
MM3 net60 B1 net36 VPW n18 W=430.00n L=180.00n
MM4 Z net60 VSS VPW n18 W=720.00n L=180.00n
MM8 net60 C1 net52 VPW n18 W=430.00n L=180.00n
MM12 net52 C2 VSS VPW n18 W=430.00n L=180.00n
MM15 net56 A2 VSS VPW n18 W=430.00n L=180.00n
MM16 net60 A1 net56 VPW n18 W=430.00n L=180.00n
.ENDS AO222UHDV1
.SUBCKT AO222UHDV2 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM1 Z net60 VDD VNW p18 W=2.02u L=180.00n
MM6 net27 A2 VDD VNW p18 W=950.0n L=180.00n
MM7 net27 A1 VDD VNW p18 W=950.0n L=180.00n
MM10 net31 B2 net27 VNW p18 W=950.0n L=180.00n
MM11 net31 B1 net27 VNW p18 W=950.0n L=180.00n
MM2 net60 C1 net31 VNW p18 W=950.0n L=180.00n
MM0 net60 C2 net31 VNW p18 W=950.0n L=180.00n
MM5 net36 B2 VSS VPW n18 W=690.00n L=180.00n
MM3 net60 B1 net36 VPW n18 W=690.00n L=180.00n
MM4 Z net60 VSS VPW n18 W=1.44u L=180.00n
MM8 net60 C1 net52 VPW n18 W=690.00n L=180.00n
MM12 net52 C2 VSS VPW n18 W=690.00n L=180.00n
MM15 net56 A2 VSS VPW n18 W=690.00n L=180.00n
MM16 net60 A1 net56 VPW n18 W=690.00n L=180.00n
.ENDS AO222UHDV2
.SUBCKT AO222UHDV3 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM1 Z net60 VDD VNW p18 W=3.03u L=180.00n
MM6 net27 A2 VDD VNW p18 W=1.01u L=180.00n
MM7 net27 A1 VDD VNW p18 W=1.01u L=180.00n
MM10 net31 B2 net27 VNW p18 W=1.01u L=180.00n
MM11 net31 B1 net27 VNW p18 W=1.01u L=180.00n
MM2 net60 C1 net31 VNW p18 W=1.01u L=180.00n
MM0 net60 C2 net31 VNW p18 W=1.01u L=180.00n
MM5 net36 B2 VSS VPW n18 W=720.00n L=180.00n
MM3 net60 B1 net36 VPW n18 W=720.00n L=180.00n
MM4 Z net60 VSS VPW n18 W=2.16u L=180.00n
MM8 net60 C1 net52 VPW n18 W=720.00n L=180.00n
MM12 net52 C2 VSS VPW n18 W=720.00n L=180.00n
MM15 net56 A2 VSS VPW n18 W=720.00n L=180.00n
MM16 net60 A1 net56 VPW n18 W=720.00n L=180.00n
.ENDS AO222UHDV3
.SUBCKT AO22UHDV0P4 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM1 Z net42 VDD VNW p18 W=490.0n L=180.00n
MM6 net25 A2 VDD VNW p18 W=490.0n L=180.00n
MM7 net25 A1 VDD VNW p18 W=490.0n L=180.00n
MM10 net42 B2 net25 VNW p18 W=490.0n L=180.00n
MM11 net42 B1 net25 VNW p18 W=490.0n L=180.00n
MM5 net30 B2 VSS VPW n18 W=0.28u L=180.00n
MM3 net42 B1 net30 VPW n18 W=0.28u L=180.00n
MM4 Z net42 VSS VPW n18 W=0.28u L=180.00n
MM15 net38 A2 VSS VPW n18 W=0.28u L=180.00n
MM16 net42 A1 net38 VPW n18 W=0.28u L=180.00n
.ENDS AO22UHDV0P4
.SUBCKT AO22UHDV0P7 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM16 net6 A1 net10 VPW n18 W=430.00n L=180.00n
MM15 net10 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 net6 B1 net18 VPW n18 W=430.00n L=180.00n
MM5 net18 B2 VSS VPW n18 W=430.00n L=180.00n
MM4 Z net6 VSS VPW n18 W=560.00n L=180.00n
MM11 net6 B1 net29 VNW p18 W=500.0n L=180.00n
MM10 net6 B2 net29 VNW p18 W=500.0n L=180.00n
MM7 net29 A1 VDD VNW p18 W=500.0n L=180.00n
MM6 net29 A2 VDD VNW p18 W=500.0n L=180.00n
MM1 Z net6 VDD VNW p18 W=790.0n L=180.00n
.ENDS AO22UHDV0P7
.SUBCKT AO22UHDV1 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM16 net6 A1 net10 VPW n18 W=430.00n L=180.00n
MM15 net10 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 net6 B1 net18 VPW n18 W=430.00n L=180.00n
MM5 net18 B2 VSS VPW n18 W=430.00n L=180.00n
MM4 Z net6 VSS VPW n18 W=720.00n L=180.00n
MM11 net6 B1 net29 VNW p18 W=580.0n L=180.00n
MM10 net6 B2 net29 VNW p18 W=580.0n L=180.00n
MM7 net29 A1 VDD VNW p18 W=580.0n L=180.00n
MM6 net29 A2 VDD VNW p18 W=580.0n L=180.00n
MM1 Z net6 VDD VNW p18 W=1.01u L=180.00n
.ENDS AO22UHDV1
.SUBCKT AO22UHDV2 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM16 net6 A1 net10 VPW n18 W=630.00n L=180.00n
MM15 net10 A2 VSS VPW n18 W=630.00n L=180.00n
MM3 net6 B1 net18 VPW n18 W=630.00n L=180.00n
MM5 net18 B2 VSS VPW n18 W=630.00n L=180.00n
MM4 Z net6 VSS VPW n18 W=1.44u L=180.00n
MM11 net6 B1 net29 VNW p18 W=950.0n L=180.00n
MM10 net6 B2 net29 VNW p18 W=950.0n L=180.00n
MM7 net29 A1 VDD VNW p18 W=950.0n L=180.00n
MM6 net29 A2 VDD VNW p18 W=950.0n L=180.00n
MM1 Z net6 VDD VNW p18 W=2.02u L=180.00n
.ENDS AO22UHDV2
.SUBCKT AO22UHDV3 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM16 net6 A1 net10 VPW n18 W=720.00n L=180.00n
MM15 net10 A2 VSS VPW n18 W=720.00n L=180.00n
MM3 net6 B1 net18 VPW n18 W=720.00n L=180.00n
MM5 net18 B2 VSS VPW n18 W=720.00n L=180.00n
MM4 Z net6 VSS VPW n18 W=2.16u L=180.00n
MM11 net6 B1 net29 VNW p18 W=1.01u L=180.00n
MM10 net6 B2 net29 VNW p18 W=1.01u L=180.00n
MM7 net29 A1 VDD VNW p18 W=1.01u L=180.00n
MM6 net29 A2 VDD VNW p18 W=1.01u L=180.00n
MM1 Z net6 VDD VNW p18 W=3.03u L=180.00n
.ENDS AO22UHDV3
.SUBCKT AO22UHDV4 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM16 net6 A1 net10 VPW n18 W=1060.00n L=180.00n
MM15 net10 A2 VSS VPW n18 W=1060.00n L=180.00n
MM3 net6 B1 net18 VPW n18 W=1060.00n L=180.00n
MM5 net18 B2 VSS VPW n18 W=1060.00n L=180.00n
MM4 Z net6 VSS VPW n18 W=2.88u L=180.00n
MM11 net6 B1 net29 VNW p18 W=1.32u L=180.00n
MM10 net6 B2 net29 VNW p18 W=1.48u L=180.00n
MM7 net29 A1 VDD VNW p18 W=1.32u L=180.00n
MM6 net29 A2 VDD VNW p18 W=1.48u L=180.00n
MM1 Z net6 VDD VNW p18 W=4.04u L=180.00n
.ENDS AO22UHDV4
.SUBCKT AO22UHDV6 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM16 net6 A1 net10 VPW n18 W=1.44u L=180.00n
MM15 net10 A2 VSS VPW n18 W=1.44u L=180.00n
MM3 net6 B1 net18 VPW n18 W=1.44u L=180.00n
MM5 net18 B2 VSS VPW n18 W=1.44u L=180.00n
MM4 Z net6 VSS VPW n18 W=4.32u L=180.00n
MM11 net6 B1 net29 VNW p18 W=2.02u L=180.00n
MM10 net6 B2 net29 VNW p18 W=2.02u L=180.00n
MM7 net29 A1 VDD VNW p18 W=2.02u L=180.00n
MM6 net29 A2 VDD VNW p18 W=2.02u L=180.00n
MM1 Z net6 VDD VNW p18 W=6.06u L=180.00n
.ENDS AO22UHDV6
.SUBCKT AO31UHDV0P4 A1 A2 A3 B Z VDD VSS VNW VPW
MM6 net10 A3 VDD VNW p18 W=490.0n L=180.00n
MM7 net38 B net10 VNW p18 W=490.0n L=180.00n
MM2 net10 A1 VDD VNW p18 W=490.0n L=180.00n
MM0 net10 A2 VDD VNW p18 W=490.0n L=180.00n
MM1 Z net38 VDD VNW p18 W=490.0n L=180.00n
MM9 net26 A3 VSS VPW n18 W=0.28u L=180.00n
MM8 net38 B VSS VPW n18 W=0.28u L=180.00n
MM5 net34 A2 net26 VPW n18 W=0.28u L=180.00n
MM3 net38 A1 net34 VPW n18 W=0.28u L=180.00n
MM4 Z net38 VSS VPW n18 W=0.28u L=180.00n
.ENDS AO31UHDV0P4
.SUBCKT AO31UHDV0P7 A1 A2 A3 B Z VDD VSS VNW VPW
MM4 Z net10 VSS VPW n18 W=560.00n L=180.00n
MM3 net10 A1 net14 VPW n18 W=430.00n L=180.00n
MM5 net14 A2 net046 VPW n18 W=430.00n L=180.00n
MM8 net10 B VSS VPW n18 W=430.00n L=180.00n
MM9 net046 A3 VSS VPW n18 W=430.00n L=180.00n
MM1 Z net10 VDD VNW p18 W=790.0n L=180.00n
MM7 net10 B net38 VNW p18 W=500.0n L=180.00n
MM0 net38 A2 VDD VNW p18 W=500.0n L=180.00n
MM2 net38 A1 VDD VNW p18 W=500.0n L=180.00n
MM6 net38 A3 VDD VNW p18 W=500.0n L=180.00n
.ENDS AO31UHDV0P7
.SUBCKT AO31UHDV1 A1 A2 A3 B Z VDD VSS VNW VPW
MM4 Z net10 VSS VPW n18 W=720.00n L=180.00n
MM3 net10 A1 net14 VPW n18 W=430.00n L=180.00n
MM5 net14 A2 net046 VPW n18 W=430.00n L=180.00n
MM8 net10 B VSS VPW n18 W=430.00n L=180.00n
MM9 net046 A3 VSS VPW n18 W=430.00n L=180.00n
MM1 Z net10 VDD VNW p18 W=1.01u L=180.00n
MM7 net10 B net38 VNW p18 W=580.0n L=180.00n
MM0 net38 A2 VDD VNW p18 W=580.0n L=180.00n
MM2 net38 A1 VDD VNW p18 W=580.0n L=180.00n
MM6 net38 A3 VDD VNW p18 W=580.0n L=180.00n
.ENDS AO31UHDV1
.SUBCKT AO31UHDV2 A1 A2 A3 B Z VDD VSS VNW VPW
MM4 Z net10 VSS VPW n18 W=1.44u L=180.00n
MM3 net10 A1 net14 VPW n18 W=630.00n L=180.00n
MM5 net14 A2 net046 VPW n18 W=630.00n L=180.00n
MM8 net10 B VSS VPW n18 W=460.00n L=180.00n
MM9 net046 A3 VSS VPW n18 W=630.00n L=180.00n
MM1 Z net10 VDD VNW p18 W=2.02u L=180.00n
MM7 net10 B net38 VNW p18 W=950.0n L=180.00n
MM0 net38 A2 VDD VNW p18 W=950.0n L=180.00n
MM2 net38 A1 VDD VNW p18 W=950.0n L=180.00n
MM6 net38 A3 VDD VNW p18 W=950.0n L=180.00n
.ENDS AO31UHDV2
.SUBCKT AO32UHDV0P7 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM11 net034 B2 VSS VPW n18 W=430.00n L=180.00n
MM10 net3 B1 net034 VPW n18 W=430.00n L=180.00n
MM9 net3 A1 net026 VPW n18 W=430.00n L=180.00n
MM8 net026 A2 net030 VPW n18 W=430.00n L=180.00n
MM7 net030 A3 VSS VPW n18 W=430.00n L=180.00n
MM0 Z net3 VSS VPW n18 W=560.00n L=180.00n
MM6 net3 B2 net054 VNW p18 W=500.00n L=180.00n
MM5 net3 B1 net054 VNW p18 W=500.00n L=180.00n
MM4 net054 A1 VDD VNW p18 W=500.00n L=180.00n
MM3 net054 A2 VDD VNW p18 W=500.00n L=180.00n
MM2 net054 A3 VDD VNW p18 W=500.00n L=180.00n
MM1 Z net3 VDD VNW p18 W=790.00n L=180.00n
.ENDS AO32UHDV0P7
.SUBCKT AO32UHDV1 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM1 Z net51 VDD VNW p18 W=1.01u L=180.00n
MM2 net19 A3 VDD VNW p18 W=580.00n L=180.00n
MM3 net19 A2 VDD VNW p18 W=580.00n L=180.00n
MM4 net19 A1 VDD VNW p18 W=580.00n L=180.00n
MM5 net51 B1 net19 VNW p18 W=580.00n L=180.00n
MM6 net51 B2 net19 VNW p18 W=580.00n L=180.00n
MM0 Z net51 VSS VPW n18 W=720.00n L=180.00n
MM10 net51 B1 net39 VPW n18 W=430.00n L=180.00n
MM11 net39 B2 VSS VPW n18 W=430.00n L=180.00n
MM7 net43 A3 VSS VPW n18 W=430.00n L=180.00n
MM8 net47 A2 net43 VPW n18 W=430.00n L=180.00n
MM9 net51 A1 net47 VPW n18 W=430.00n L=180.00n
.ENDS AO32UHDV1
.SUBCKT AO32UHDV2 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM9 net7 A1 net11 VPW n18 W=630.00n L=180.00n
MM8 net11 A2 net15 VPW n18 W=630.00n L=180.00n
MM7 net15 A3 VSS VPW n18 W=630.00n L=180.00n
MM11 net19 B2 VSS VPW n18 W=630.00n L=180.00n
MM10 net7 B1 net19 VPW n18 W=630.00n L=180.00n
MM0 Z net7 VSS VPW n18 W=1.44u L=180.00n
MM6 net7 B2 net39 VNW p18 W=950.00n L=180.00n
MM5 net7 B1 net39 VNW p18 W=950.00n L=180.00n
MM4 net39 A1 VDD VNW p18 W=950.00n L=180.00n
MM3 net39 A2 VDD VNW p18 W=950.00n L=180.00n
MM2 net39 A3 VDD VNW p18 W=950.00n L=180.00n
MM1 Z net7 VDD VNW p18 W=2.02u L=180.00n
.ENDS AO32UHDV2
.SUBCKT AO32UHDV3 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM1 Z net51 VDD VNW p18 W=3.03u L=180.00n
MM2 net19 A3 VDD VNW p18 W=1.01u L=180.00n
MM3 net19 A2 VDD VNW p18 W=1.01u L=180.00n
MM4 net19 A1 VDD VNW p18 W=1.01u L=180.00n
MM5 net51 B1 net19 VNW p18 W=1.01u L=180.00n
MM6 net51 B2 net19 VNW p18 W=1.01u L=180.00n
MM0 Z net51 VSS VPW n18 W=2.16u L=180.00n
MM10 net51 B1 net39 VPW n18 W=720.00n L=180.00n
MM11 net39 B2 VSS VPW n18 W=720.00n L=180.00n
MM7 net43 A3 VSS VPW n18 W=720.00n L=180.00n
MM8 net47 A2 net43 VPW n18 W=720.00n L=180.00n
MM9 net51 A1 net47 VPW n18 W=720.00n L=180.00n
.ENDS AO32UHDV3
.SUBCKT AO32UHDV4 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM9 net7 A1 net11 VPW n18 W=1060.0n L=180.00n
MM8 net11 A2 net15 VPW n18 W=1060.0n L=180.00n
MM7 net15 A3 VSS VPW n18 W=1060.0n L=180.00n
MM11 net19 B2 VSS VPW n18 W=1060.0n L=180.00n
MM10 net7 B1 net19 VPW n18 W=1060.0n L=180.00n
MM0 Z net7 VSS VPW n18 W=2.88u L=180.00n
MM6 net7 B2 net39 VNW p18 W=1.82u L=180.00n
MM5 net7 B1 net39 VNW p18 W=1.82u L=180.00n
MM4 net39 A1 VDD VNW p18 W=1.49u L=180.00n
MM3 net39 A2 VDD VNW p18 W=1.49u L=180.00n
MM2 net39 A3 VDD VNW p18 W=1.49u L=180.00n
MM1 Z net7 VDD VNW p18 W=4.04u L=180.00n
.ENDS AO32UHDV4
.SUBCKT AO33UHDV0P7 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM12 net60 B3 net24 VNW p18 W=500.00n L=180.00n
MM1 Z net60 VDD VNW p18 W=790.00n L=180.00n
MM2 net24 A3 VDD VNW p18 W=500.00n L=180.00n
MM3 net24 A2 VDD VNW p18 W=500.00n L=180.00n
MM4 net24 A1 VDD VNW p18 W=500.00n L=180.00n
MM5 net60 B1 net24 VNW p18 W=500.00n L=180.00n
MM6 net60 B2 net24 VNW p18 W=500.00n L=180.00n
MM0 Z net60 VSS VPW n18 W=560.00n L=180.00n
MM10 net60 B1 net40 VPW n18 W=430.00n L=180.00n
MM11 net40 B2 net44 VPW n18 W=430.00n L=180.00n
MM7 net52 A3 VSS VPW n18 W=430.00n L=180.00n
MM8 net56 A2 net52 VPW n18 W=430.00n L=180.00n
MM9 net60 A1 net56 VPW n18 W=430.00n L=180.00n
MM13 net44 B3 VSS VPW n18 W=430.00n L=180.00n
.ENDS AO33UHDV0P7
.SUBCKT AO33UHDV1 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM9 net8 A1 net12 VPW n18 W=430.00n L=180.00n
MM8 net12 A2 net16 VPW n18 W=430.00n L=180.00n
MM7 net16 A3 VSS VPW n18 W=430.00n L=180.00n
MM0 Z net8 VSS VPW n18 W=720.0n L=180.00n
MM13 net24 B3 VSS VPW n18 W=430.00n L=180.00n
MM11 net28 B2 net24 VPW n18 W=430.00n L=180.00n
MM10 net8 B1 net28 VPW n18 W=430.00n L=180.00n
MM6 net8 B2 net44 VNW p18 W=580.00n L=180.00n
MM5 net8 B1 net44 VNW p18 W=580.00n L=180.00n
MM4 net44 A1 VDD VNW p18 W=580.00n L=180.00n
MM3 net44 A2 VDD VNW p18 W=580.00n L=180.00n
MM2 net44 A3 VDD VNW p18 W=580.00n L=180.00n
MM1 Z net8 VDD VNW p18 W=1.01u L=180.00n
MM12 net8 B3 net44 VNW p18 W=580.00n L=180.00n
.ENDS AO33UHDV1
.SUBCKT AO33UHDV2 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM12 net60 B3 net24 VNW p18 W=950.00n L=180.00n
MM1 Z net60 VDD VNW p18 W=2.02u L=180.00n
MM2 net24 A3 VDD VNW p18 W=950.00n L=180.00n
MM3 net24 A2 VDD VNW p18 W=950.00n L=180.00n
MM4 net24 A1 VDD VNW p18 W=950.00n L=180.00n
MM5 net60 B1 net24 VNW p18 W=950.00n L=180.00n
MM6 net60 B2 net24 VNW p18 W=950.00n L=180.00n
MM10 net60 B1 net40 VPW n18 W=630.00n L=180.00n
MM11 net40 B2 net44 VPW n18 W=630.00n L=180.00n
MM13 net44 B3 VSS VPW n18 W=630.00n L=180.00n
MM0 Z net60 VSS VPW n18 W=1.44u L=180.00n
MM7 net52 A3 VSS VPW n18 W=630.00n L=180.00n
MM8 net56 A2 net52 VPW n18 W=630.00n L=180.00n
MM9 net60 A1 net56 VPW n18 W=630.00n L=180.00n
.ENDS AO33UHDV2
.SUBCKT AO33UHDV3 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM9 net8 A1 net12 VPW n18 W=720.00n L=180.00n
MM8 net12 A2 net16 VPW n18 W=720.00n L=180.00n
MM7 net16 A3 VSS VPW n18 W=720.00n L=180.00n
MM0 Z net8 VSS VPW n18 W=2.16u L=180.00n
MM13 net24 B3 VSS VPW n18 W=720.00n L=180.00n
MM11 net28 B2 net24 VPW n18 W=720.00n L=180.00n
MM10 net8 B1 net28 VPW n18 W=720.00n L=180.00n
MM6 net8 B2 net44 VNW p18 W=1.01u L=180.00n
MM5 net8 B1 net44 VNW p18 W=1.01u L=180.00n
MM4 net44 A1 VDD VNW p18 W=1.01u L=180.00n
MM3 net44 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net44 A3 VDD VNW p18 W=1.01u L=180.00n
MM1 Z net8 VDD VNW p18 W=3.03u L=180.00n
MM12 net8 B3 net44 VNW p18 W=1.01u L=180.00n
.ENDS AO33UHDV3
.SUBCKT AO33UHDV4 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM12 net60 B3 net24 VNW p18 W=1.49u L=180.00n
MM1 Z net60 VDD VNW p18 W=4.04u L=180.00n
MM2 net24 A3 VDD VNW p18 W=1.49u L=180.00n
MM3 net24 A2 VDD VNW p18 W=1.49u L=180.00n
MM4 net24 A1 VDD VNW p18 W=1.49u L=180.00n
MM5 net60 B1 net24 VNW p18 W=1.49u L=180.00n
MM6 net60 B2 net24 VNW p18 W=1.49u L=180.00n
MM10 net60 B1 net40 VPW n18 W=1060.00n L=180.00n
MM11 net40 B2 net44 VPW n18 W=1060.00n L=180.00n
MM13 net44 B3 VSS VPW n18 W=1060.00n L=180.00n
MM0 Z net60 VSS VPW n18 W=2.88u L=180.00n
MM7 net52 A3 VSS VPW n18 W=1060.00n L=180.00n
MM8 net56 A2 net52 VPW n18 W=1060.00n L=180.00n
MM9 net60 A1 net56 VPW n18 W=1060.00n L=180.00n
.ENDS AO33UHDV4
.SUBCKT AOI211UHDV0P4 A1 A2 B C ZN VDD VSS VNW VPW
MM3 ZN A1 net10 VPW n18 W=0.28u L=180.00n
MM5 net10 A2 VSS VPW n18 W=0.28u L=180.00n
MM8 ZN B VSS VPW n18 W=0.28u L=180.00n
MM9 ZN C VSS VPW n18 W=0.28u L=180.00n
MM0 net26 A2 VDD VNW p18 W=490.0n L=180.00n
MM2 net26 A1 VDD VNW p18 W=490.0n L=180.00n
MM6 net37 B net26 VNW p18 W=490.0n L=180.00n
MM7 ZN C net37 VNW p18 W=490.0n L=180.00n
.ENDS AOI211UHDV0P4
.SUBCKT AOI211UHDV0P7 A1 A2 B C ZN VDD VSS VNW VPW
MM7 ZN C net9 VNW p18 W=760.0n L=180.00n
MM6 net9 B net14 VNW p18 W=760.0n L=180.00n
MM2 net14 A1 VDD VNW p18 W=760.0n L=180.00n
MM0 net14 A2 VDD VNW p18 W=760.0n L=180.00n
MM9 ZN C VSS VPW n18 W=500.00n L=180.00n
MM8 ZN B VSS VPW n18 W=500.00n L=180.00n
MM5 net30 A2 VSS VPW n18 W=500.00n L=180.00n
MM3 ZN A1 net30 VPW n18 W=500.00n L=180.00n
.ENDS AOI211UHDV0P7
.SUBCKT AOI211UHDV1 A1 A2 B C ZN VDD VSS VNW VPW
MM3 ZN A1 net10 VPW n18 W=720.00n L=180.00n
MM5 net10 A2 VSS VPW n18 W=720.00n L=180.00n
MM8 ZN B VSS VPW n18 W=720.00n L=180.00n
MM9 ZN C VSS VPW n18 W=720.00n L=180.00n
MM0 net26 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net26 A1 VDD VNW p18 W=1.01u L=180.00n
MM6 net37 B net26 VNW p18 W=1.01u L=180.00n
MM7 ZN C net37 VNW p18 W=1.01u L=180.00n
.ENDS AOI211UHDV1
.SUBCKT AOI211UHDV2 A1 A2 B C ZN VDD VSS VNW VPW
MM3 ZN A1 net10 VPW n18 W=1.44u L=180.00n
MM5 net10 A2 VSS VPW n18 W=1.44u L=180.00n
MM8 ZN B VSS VPW n18 W=1.44u L=180.00n
MM9 ZN C VSS VPW n18 W=1.44u L=180.00n
MM0 net26 A2 VDD VNW p18 W=2.02u L=180.00n
MM2 net26 A1 VDD VNW p18 W=2.02u L=180.00n
MM6 net37 B net26 VNW p18 W=2.02u L=180.00n
MM7 ZN C net37 VNW p18 W=1.95u L=180.00n
.ENDS AOI211UHDV2
.SUBCKT AOI211UHDV3 A1 A2 B C ZN VDD VSS VNW VPW
MM3 ZN A1 net10 VPW n18 W=2.16u L=180.00n
MM5 net10 A2 VSS VPW n18 W=2.16u L=180.00n
MM8 ZN B VSS VPW n18 W=2.16u L=180.00n
MM9 ZN C VSS VPW n18 W=2.16u L=180.00n
MM0 net26 A2 VDD VNW p18 W=3.03u L=180.00n
MM2 net26 A1 VDD VNW p18 W=2.96u L=180.00n
MM6 net37 B net26 VNW p18 W=3.03u L=180.00n
MM7 ZN C net37 VNW p18 W=2.96u L=180.00n
.ENDS AOI211UHDV3
.SUBCKT AOI21BUHDV0P4 A B1 B2 ZN VDD VSS VNW VPW
MM3 ZN B1 net9 VPW n18 W=0.28u L=180.00n
MM5 net9 B2 VSS VPW n18 W=0.28u L=180.00n
MM8 ZN net17 VSS VPW n18 W=0.28u L=180.00n
MM6 net17 A VSS VPW n18 W=0.28u L=180.00n
MM1 ZN net17 net29 VNW p18 W=0.5u L=180.00n
MM0 net29 B2 VDD VNW p18 W=0.5u L=180.00n
MM2 net29 B1 VDD VNW p18 W=0.5u L=180.00n
MM4 net17 A VDD VNW p18 W=0.49u L=180.00n
.ENDS AOI21BUHDV0P4
.SUBCKT AOI21BUHDV0P7 A B1 B2 ZN VDD VSS VNW VPW
MM3 ZN B1 net9 VPW n18 W=0.44u L=180.00n
MM5 net9 B2 VSS VPW n18 W=0.44u L=180.00n
MM8 ZN net17 VSS VPW n18 W=560.00n L=180.00n
MM6 net17 A VSS VPW n18 W=0.42u L=180.00n
MM1 ZN net17 net29 VNW p18 W=780.00n L=180.00n
MM0 net29 B2 VDD VNW p18 W=670.00n L=180.00n
MM2 net29 B1 VDD VNW p18 W=670.00n L=180.00n
MM4 net17 A VDD VNW p18 W=0.515u L=180.00n
.ENDS AOI21BUHDV0P7
.SUBCKT AOI21BUHDV1 A B1 B2 ZN VDD VSS VNW VPW
MM3 ZN B1 net9 VPW n18 W=720.00n L=180.00n
MM5 net9 B2 VSS VPW n18 W=720.00n L=180.00n
MM8 ZN net17 VSS VPW n18 W=720.00n L=180.00n
MM6 net17 A VSS VPW n18 W=430.00n L=180.00n
MM1 ZN net17 net29 VNW p18 W=1.01u L=180.00n
MM0 net29 B2 VDD VNW p18 W=1.01u L=180.00n
MM2 net29 B1 VDD VNW p18 W=1.01u L=180.00n
MM4 net17 A VDD VNW p18 W=0.59u L=180.00n
.ENDS AOI21BUHDV1
.SUBCKT AOI21BUHDV2 A B1 B2 ZN VDD VSS VNW VPW
MM4 net21 A VDD VNW p18 W=0.965u L=180.00n
MM2 net9 B1 VDD VNW p18 W=1.89u L=180.00n
MM0 net9 B2 VDD VNW p18 W=2.01u L=180.00n
MM1 ZN net21 net9 VNW p18 W=2.01u L=180.00n
MM6 net21 A VSS VPW n18 W=630.00n L=180.00n
MM8 ZN net21 VSS VPW n18 W=1.44u L=180.00n
MM5 net29 B2 VSS VPW n18 W=1.44u L=180.00n
MM3 ZN B1 net29 VPW n18 W=1.44u L=180.00n
.ENDS AOI21BUHDV2
.SUBCKT AOI21UHDV0P4 A1 A2 B ZN VDD VSS VNW VPW
MM1 ZN B net4 VNW p18 W=0.475u L=180.00n
MM2 net4 A1 VDD VNW p18 W=0.475u L=180.00n
MM0 net4 A2 VDD VNW p18 W=0.475u L=180.00n
MM8 ZN B VSS VPW n18 W=0.28u L=180.00n
MM5 net20 A2 VSS VPW n18 W=0.28u L=180.00n
MM3 ZN A1 net20 VPW n18 W=0.28u L=180.00n
.ENDS AOI21UHDV0P4
.SUBCKT AOI21UHDV0P7 A1 A2 B ZN VDD VSS VNW VPW
MM3 ZN A1 net8 VPW n18 W=560.00n L=180.00n
MM5 net8 A2 VSS VPW n18 W=560.00n L=180.00n
MM8 ZN B VSS VPW n18 W=560.00n L=180.00n
MM1 ZN B net24 VNW p18 W=675.00n L=180.00n
MM0 net24 A2 VDD VNW p18 W=0.475u L=180.00n
MM2 net24 A1 VDD VNW p18 W=675.00n L=180.00n
.ENDS AOI21UHDV0P7
.SUBCKT AOI21UHDV1 A1 A2 B ZN VDD VSS VNW VPW
MM3 ZN A1 net8 VPW n18 W=720.00n L=180.00n
MM5 net8 A2 VSS VPW n18 W=720.00n L=180.00n
MM8 ZN B VSS VPW n18 W=720.00n L=180.00n
MM1 ZN B net24 VNW p18 W=1.01u L=180.00n
MM0 net24 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net24 A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS AOI21UHDV1
.SUBCKT AOI21UHDV2 A1 A2 B ZN VDD VSS VNW VPW
MM3 ZN A1 net8 VPW n18 W=1.44u L=180.00n
MM5 net8 A2 VSS VPW n18 W=1.44u L=180.00n
MM8 ZN B VSS VPW n18 W=1.44u L=180.00n
MM1 ZN B net24 VNW p18 W=2.02u L=180.00n
MM0 net24 A2 VDD VNW p18 W=2.02u L=180.00n
MM2 net24 A1 VDD VNW p18 W=2.02u L=180.00n
.ENDS AOI21UHDV2
.SUBCKT AOI21UHDV3 A1 A2 B ZN VDD VSS VNW VPW
MM3 ZN A1 net8 VPW n18 W=2.11u L=180.00n
MM5 net8 A2 VSS VPW n18 W=2.11u L=180.00n
MM8 ZN B VSS VPW n18 W=2.085u L=180.00n
MM1 ZN B net24 VNW p18 W=3.03u L=180.00n
MM0 net24 A2 VDD VNW p18 W=2.96u L=180.00n
MM2 net24 A1 VDD VNW p18 W=3.03u L=180.00n
.ENDS AOI21UHDV3
.SUBCKT AOI21UHDV4 A1 A2 B ZN VDD VSS VNW VPW
MM3 ZN A1 net8 VPW n18 W=2.88u L=180.00n
MM5 net8 A2 VSS VPW n18 W=2.88u L=180.00n
MM8 ZN B VSS VPW n18 W=2.88u L=180.00n
MM1 ZN B net24 VNW p18 W=4.04u L=180.00n
MM0 net24 A2 VDD VNW p18 W=3.97u L=180.00n
MM2 net24 A1 VDD VNW p18 W=4.04u L=180.00n
.ENDS AOI21UHDV4
.SUBCKT AOI21UHDV6 A1 A2 B ZN VDD VSS VNW VPW
MM3 ZN A1 net8 VPW n18 W=4.32u L=180.00n
MM5 net8 A2 VSS VPW n18 W=4.32u L=180.00n
MM8 ZN B VSS VPW n18 W=4.32u L=180.00n
MM1 ZN B net24 VNW p18 W=6.06u L=180.00n
MM0 net24 A2 VDD VNW p18 W=5.92u L=180.00n
MM2 net24 A1 VDD VNW p18 W=6.06u L=180.00n
.ENDS AOI21UHDV6
.SUBCKT AOI221UHDV0P4 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM3 ZN A1 net15 VPW n18 W=0.28u L=180.00n
MM5 net15 A2 VSS VPW n18 W=0.28u L=180.00n
MM8 ZN B1 net7 VPW n18 W=0.28u L=180.00n
MM9 ZN C VSS VPW n18 W=0.28u L=180.00n
MM6 net7 B2 VSS VPW n18 W=0.28u L=180.00n
MM0 net30 A2 VDD VNW p18 W=490.0n L=180.00n
MM2 net30 A1 VDD VNW p18 W=490.0n L=180.00n
MM1 net27 B2 net30 VNW p18 W=490.0n L=180.00n
MM7 ZN C net27 VNW p18 W=490.0n L=180.00n
MM4 net27 B1 net30 VNW p18 W=490.0n L=180.00n
.ENDS AOI221UHDV0P4
.SUBCKT AOI221UHDV0P7 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM7 ZN C net23 VNW p18 W=675.00n L=180.00n
MM2 net26 A1 VDD VNW p18 W=0.675u L=180.00n
MM0 net26 A2 VDD VNW p18 W=0.675u L=180.00n
MM1 net23 B2 net26 VNW p18 W=0.675u L=180.00n
MM4 net23 B1 net26 VNW p18 W=0.675u L=180.00n
MM9 ZN C VSS VPW n18 W=560.00n L=180.00n
MM8 ZN B1 net43 VPW n18 W=560.00n L=180.00n
MM5 net35 A2 VSS VPW n18 W=560.00n L=180.00n
MM3 ZN A1 net35 VPW n18 W=560.00n L=180.00n
MM6 net43 B2 VSS VPW n18 W=560.00n L=180.00n
.ENDS AOI221UHDV0P7
.SUBCKT AOI221UHDV1 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM6 net7 B2 VSS VPW n18 W=720.00n L=180.00n
MM3 ZN A1 net15 VPW n18 W=720.00n L=180.00n
MM5 net15 A2 VSS VPW n18 W=720.00n L=180.00n
MM8 ZN B1 net7 VPW n18 W=720.00n L=180.00n
MM9 ZN C VSS VPW n18 W=720.00n L=180.00n
MM4 net27 B1 net30 VNW p18 W=1.01u L=180.00n
MM1 net27 B2 net30 VNW p18 W=1.01u L=180.00n
MM0 net30 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net30 A1 VDD VNW p18 W=1.01u L=180.00n
MM7 ZN C net27 VNW p18 W=1.01u L=180.00n
.ENDS AOI221UHDV1
.SUBCKT AOI221UHDV2 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM6 net7 B2 VSS VPW n18 W=1.44u L=180.00n
MM3 ZN A1 net15 VPW n18 W=1.44u L=180.00n
MM5 net15 A2 VSS VPW n18 W=1.44u L=180.00n
MM8 ZN B1 net7 VPW n18 W=1.44u L=180.00n
MM9 ZN C VSS VPW n18 W=1.44u L=180.00n
MM4 net27 B1 net30 VNW p18 W=2.02u L=180.00n
MM1 net27 B2 net30 VNW p18 W=2.02u L=180.00n
MM0 net30 A2 VDD VNW p18 W=2.02u L=180.00n
MM2 net30 A1 VDD VNW p18 W=2.02u L=180.00n
MM7 ZN C net27 VNW p18 W=2.02u L=180.00n
.ENDS AOI221UHDV2
.SUBCKT AOI221UHDV3 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM6 net7 B2 VSS VPW n18 W=2.16u L=180.00n
MM3 ZN A1 net15 VPW n18 W=2.16u L=180.00n
MM5 net15 A2 VSS VPW n18 W=2.16u L=180.00n
MM8 ZN B1 net7 VPW n18 W=2.16u L=180.00n
MM9 ZN C VSS VPW n18 W=2.14u L=180.00n
MM4 net27 B1 net30 VNW p18 W=3.03u L=180.00n
MM1 net27 B2 net30 VNW p18 W=2.96u L=180.00n
MM0 net30 A2 VDD VNW p18 W=3.03u L=180.00n
MM2 net30 A1 VDD VNW p18 W=3.03u L=180.00n
MM7 ZN C net27 VNW p18 W=3.03u L=180.00n
.ENDS AOI221UHDV3
.SUBCKT AOI221UHDV4 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM6 net7 B2 VSS VPW n18 W=2.88u L=180.00n
MM3 ZN A1 net15 VPW n18 W=2.88u L=180.00n
MM5 net15 A2 VSS VPW n18 W=2.88u L=180.00n
MM8 ZN B1 net7 VPW n18 W=2.88u L=180.00n
MM9 ZN C VSS VPW n18 W=2.88u L=180.00n
MM4 net27 B1 net30 VNW p18 W=4.04u L=180.00n
MM1 net27 B2 net30 VNW p18 W=3.97u L=180.00n
MM0 net30 A2 VDD VNW p18 W=4.03u L=180.00n
MM2 net30 A1 VDD VNW p18 W=4.04u L=180.00n
MM7 ZN C net27 VNW p18 W=4.11u L=180.00n
.ENDS AOI221UHDV4
.SUBCKT AOI222UHDV0P4 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM10 net19 B2 net31 VNW p18 W=490.0n L=180.00n
MM7 net31 C1 VDD VNW p18 W=490.0n L=180.00n
MM2 ZN A1 net19 VNW p18 W=490.0n L=180.00n
MM0 ZN A2 net19 VNW p18 W=490.0n L=180.00n
MM6 net31 C2 VDD VNW p18 W=490.0n L=180.00n
MM11 net19 B1 net31 VNW p18 W=490.0n L=180.00n
MM12 net32 A2 VSS VPW n18 W=0.28u L=180.00n
MM8 ZN A1 net32 VPW n18 W=0.28u L=180.00n
MM5 net40 B2 VSS VPW n18 W=0.28u L=180.00n
MM3 ZN B1 net40 VPW n18 W=0.28u L=180.00n
MM15 net48 C2 VSS VPW n18 W=0.28u L=180.00n
MM16 ZN C1 net48 VPW n18 W=0.28u L=180.00n
.ENDS AOI222UHDV0P4
.SUBCKT AOI222UHDV0P7 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM16 ZN C1 net12 VPW n18 W=0.475u L=180.00n
MM15 net12 C2 VSS VPW n18 W=0.475u L=180.00n
MM3 ZN B1 net20 VPW n18 W=0.475u L=180.00n
MM5 net20 B2 VSS VPW n18 W=0.475u L=180.00n
MM8 ZN A1 net28 VPW n18 W=0.475u L=180.00n
MM12 net28 A2 VSS VPW n18 W=0.475u L=180.00n
MM11 net47 B1 net35 VNW p18 W=0.475u L=180.00n
MM6 net35 C2 VDD VNW p18 W=675.00n L=180.00n
MM0 ZN A2 net47 VNW p18 W=0.475u L=180.00n
MM2 ZN A1 net47 VNW p18 W=0.475u L=180.00n
MM7 net35 C1 VDD VNW p18 W=675.00n L=180.00n
MM10 net47 B2 net35 VNW p18 W=0.475u L=180.00n
.ENDS AOI222UHDV0P7
.SUBCKT AOI222UHDV1 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM16 ZN C1 net12 VPW n18 W=720.00n L=180.00n
MM15 net12 C2 VSS VPW n18 W=720.00n L=180.00n
MM3 ZN B1 net20 VPW n18 W=720.00n L=180.00n
MM5 net20 B2 VSS VPW n18 W=720.00n L=180.00n
MM8 ZN A1 net28 VPW n18 W=720.00n L=180.00n
MM12 net28 A2 VSS VPW n18 W=720.00n L=180.00n
MM11 net47 B1 net35 VNW p18 W=1.01u L=180.00n
MM6 net35 C2 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN A2 net47 VNW p18 W=1.01u L=180.00n
MM2 ZN A1 net47 VNW p18 W=1.01u L=180.00n
MM7 net35 C1 VDD VNW p18 W=1.01u L=180.00n
MM10 net47 B2 net35 VNW p18 W=1.01u L=180.00n
.ENDS AOI222UHDV1
.SUBCKT AOI222UHDV2 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM16 ZN C1 net12 VPW n18 W=1.44u L=180.00n
MM15 net12 C2 VSS VPW n18 W=1.44u L=180.00n
MM3 ZN B1 net20 VPW n18 W=1.44u L=180.00n
MM5 net20 B2 VSS VPW n18 W=1.44u L=180.00n
MM8 ZN A1 net28 VPW n18 W=1.44u L=180.00n
MM12 net28 A2 VSS VPW n18 W=1.44u L=180.00n
MM11 net47 B1 net35 VNW p18 W=2.02u L=180.00n
MM6 net35 C2 VDD VNW p18 W=2.02u L=180.00n
MM0 ZN A2 net47 VNW p18 W=2.02u L=180.00n
MM2 ZN A1 net47 VNW p18 W=2.02u L=180.00n
MM7 net35 C1 VDD VNW p18 W=2.02u L=180.00n
MM10 net47 B2 net35 VNW p18 W=2.02u L=180.00n
.ENDS AOI222UHDV2
.SUBCKT AOI222UHDV3 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM16 ZN C1 net12 VPW n18 W=2.16u L=180.00n
MM15 net12 C2 VSS VPW n18 W=2.16u L=180.00n
MM3 ZN B1 net20 VPW n18 W=2.16u L=180.00n
MM5 net20 B2 VSS VPW n18 W=2.16u L=180.00n
MM8 ZN A1 net28 VPW n18 W=2.16u L=180.00n
MM12 net28 A2 VSS VPW n18 W=2.16u L=180.00n
MM11 net47 B1 net35 VNW p18 W=2.995u L=180.00n
MM6 net35 C2 VDD VNW p18 W=3.03u L=180.00n
MM0 ZN A2 net47 VNW p18 W=2.96u L=180.00n
MM2 ZN A1 net47 VNW p18 W=3.03u L=180.00n
MM7 net35 C1 VDD VNW p18 W=2.96u L=180.00n
MM10 net47 B2 net35 VNW p18 W=2.96u L=180.00n
.ENDS AOI222UHDV3
.SUBCKT AOI22BBUHDV0P4 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM10 ZN B1 net95 VNW p18 W=490.0n L=180.00n
MM5 net95 net120 VDD VNW p18 W=490.0n L=180.00n
MM3 ZN B2 net95 VNW p18 W=490.0n L=180.00n
MM1 net120 A1 net103 VNW p18 W=490.0n L=180.00n
MM4 net103 A2 VDD VNW p18 W=490.0n L=180.00n
MM9 ZN net120 VSS VPW n18 W=0.28u L=180.00n
MM2 net104 B2 VSS VPW n18 W=0.28u L=180.00n
MM0 ZN B1 net104 VPW n18 W=0.28u L=180.00n
MM8 net120 A1 VSS VPW n18 W=0.28u L=180.00n
MM6 net120 A2 VSS VPW n18 W=0.28u L=180.00n
.ENDS AOI22BBUHDV0P4
.SUBCKT AOI22BBUHDV0P7 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM8 net6 A1 VSS VPW n18 W=430.00n L=180.00n
MM6 net6 A2 VSS VPW n18 W=430.00n L=180.00n
MM9 ZN net6 VSS VPW n18 W=560.00n L=180.00n
MM0 ZN B1 net22 VPW n18 W=560.00n L=180.00n
MM2 net22 B2 VSS VPW n18 W=560.00n L=180.00n
MM1 net6 A1 net29 VNW p18 W=500.0n L=180.00n
MM4 net29 A2 VDD VNW p18 W=500.0n L=180.00n
MM3 ZN B2 net37 VNW p18 W=790.0n L=180.00n
MM10 ZN B1 net37 VNW p18 W=790.0n L=180.00n
MM5 net37 net6 VDD VNW p18 W=790.0n L=180.00n
.ENDS AOI22BBUHDV0P7
.SUBCKT AOI22BBUHDV1 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM8 net6 A1 VSS VPW n18 W=430.00n L=180.00n
MM6 net6 A2 VSS VPW n18 W=430.00n L=180.00n
MM9 ZN net6 VSS VPW n18 W=720.00n L=180.00n
MM0 ZN B1 net22 VPW n18 W=720.00n L=180.00n
MM2 net22 B2 VSS VPW n18 W=720.00n L=180.00n
MM1 net6 A1 net29 VNW p18 W=580.0n L=180.00n
MM4 net29 A2 VDD VNW p18 W=580.0n L=180.00n
MM3 ZN B2 net37 VNW p18 W=1.01u L=180.00n
MM10 ZN B1 net37 VNW p18 W=1.01u L=180.00n
MM5 net37 net6 VDD VNW p18 W=1.01u L=180.00n
.ENDS AOI22BBUHDV1
.SUBCKT AOI22BBUHDV2 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM8 net6 A1 VSS VPW n18 W=630.00n L=180.00n
MM6 net6 A2 VSS VPW n18 W=630.00n L=180.00n
MM9 ZN net6 VSS VPW n18 W=1.44u L=180.00n
MM0 ZN B1 net22 VPW n18 W=1.5u L=180.00n
MM2 net22 B2 VSS VPW n18 W=1.44u L=180.00n
MM1 net6 A1 net29 VNW p18 W=950.0n L=180.00n
MM4 net29 A2 VDD VNW p18 W=950.0n L=180.00n
MM3 ZN B2 net37 VNW p18 W=1.89u L=180.00n
MM10 ZN B1 net37 VNW p18 W=1.89u L=180.00n
MM5 net37 net6 VDD VNW p18 W=2.01u L=180.00n
.ENDS AOI22BBUHDV2
.SUBCKT AOI22UHDV0P4 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM16 ZN A1 net10 VPW n18 W=0.28u L=180.00n
MM15 net10 A2 VSS VPW n18 W=0.28u L=180.00n
MM3 ZN B1 net18 VPW n18 W=0.28u L=180.00n
MM5 net18 B2 VSS VPW n18 W=0.28u L=180.00n
MM11 ZN B1 net25 VNW p18 W=490.0n L=180.00n
MM10 ZN B2 net25 VNW p18 W=490.0n L=180.00n
MM7 net25 A1 VDD VNW p18 W=490.0n L=180.00n
MM6 net25 A2 VDD VNW p18 W=490.0n L=180.00n
.ENDS AOI22UHDV0P4
.SUBCKT AOI22UHDV0P7 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM6 net21 A2 VDD VNW p18 W=0.675u L=180.00n
MM7 net21 A1 VDD VNW p18 W=0.675u L=180.00n
MM10 ZN B2 net21 VNW p18 W=0.675u L=180.00n
MM11 ZN B1 net21 VNW p18 W=0.675u L=180.00n
MM5 net22 B2 VSS VPW n18 W=560.00n L=180.00n
MM3 ZN B1 net22 VPW n18 W=560.00n L=180.00n
MM15 net30 A2 VSS VPW n18 W=560.00n L=180.00n
MM16 ZN A1 net30 VPW n18 W=560.00n L=180.00n
.ENDS AOI22UHDV0P7
.SUBCKT AOI22UHDV1 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM6 net21 A2 VDD VNW p18 W=1.01u L=180.00n
MM7 net21 A1 VDD VNW p18 W=1.01u L=180.00n
MM10 ZN B2 net21 VNW p18 W=1.01u L=180.00n
MM11 ZN B1 net21 VNW p18 W=1.01u L=180.00n
MM5 net22 B2 VSS VPW n18 W=720.00n L=180.00n
MM3 ZN B1 net22 VPW n18 W=720.00n L=180.00n
MM15 net30 A2 VSS VPW n18 W=720.00n L=180.00n
MM16 ZN A1 net30 VPW n18 W=720.00n L=180.00n
.ENDS AOI22UHDV1
.SUBCKT AOI22UHDV2 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM6 net21 A2 VDD VNW p18 W=2.02u L=180.00n
MM7 net21 A1 VDD VNW p18 W=2.02u L=180.00n
MM10 ZN B2 net21 VNW p18 W=2.02u L=180.00n
MM11 ZN B1 net21 VNW p18 W=2.02u L=180.00n
MM5 net22 B2 VSS VPW n18 W=1.44u L=180.00n
MM3 ZN B1 net22 VPW n18 W=1.44u L=180.00n
MM15 net30 A2 VSS VPW n18 W=1.44u L=180.00n
MM16 ZN A1 net30 VPW n18 W=1.44u L=180.00n
.ENDS AOI22UHDV2
.SUBCKT AOI22UHDV3 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM6 net21 A2 VDD VNW p18 W=3.03u L=180.00n
MM7 net21 A1 VDD VNW p18 W=3.03u L=180.00n
MM10 ZN B2 net21 VNW p18 W=2.96u L=180.00n
MM11 ZN B1 net21 VNW p18 W=3.03u L=180.00n
MM5 net22 B2 VSS VPW n18 W=2.16u L=180.00n
MM3 ZN B1 net22 VPW n18 W=2.16u L=180.00n
MM15 net30 A2 VSS VPW n18 W=2.16u L=180.00n
MM16 ZN A1 net30 VPW n18 W=2.16u L=180.00n
.ENDS AOI22UHDV3
.SUBCKT AOI22UHDV4 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM6 net21 A2 VDD VNW p18 W=4.03u L=180.00n
MM7 net21 A1 VDD VNW p18 W=4.04u L=180.00n
MM10 ZN B2 net21 VNW p18 W=3.97u L=180.00n
MM11 ZN B1 net21 VNW p18 W=4.04u L=180.00n
MM5 net22 B2 VSS VPW n18 W=2.88u L=180.00n
MM3 ZN B1 net22 VPW n18 W=2.88u L=180.00n
MM15 net30 A2 VSS VPW n18 W=2.88u L=180.00n
MM16 ZN A1 net30 VPW n18 W=2.88u L=180.00n
.ENDS AOI22UHDV4
.SUBCKT AOI22UHDV6 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM6 net21 A2 VDD VNW p18 W=6.06u L=180.00n
MM7 net21 A1 VDD VNW p18 W=6.06u L=180.00n
MM10 ZN B2 net21 VNW p18 W=5.92u L=180.00n
MM11 ZN B1 net21 VNW p18 W=6.025u L=180.00n
MM5 net22 B2 VSS VPW n18 W=4.32u L=180.00n
MM3 ZN B1 net22 VPW n18 W=4.32u L=180.00n
MM15 net30 A2 VSS VPW n18 W=4.32u L=180.00n
MM16 ZN A1 net30 VPW n18 W=4.32u L=180.00n
.ENDS AOI22UHDV6
.SUBCKT AOI22XBUHDV0P4 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM5 ZN B1 net9 VNW p18 W=475.00n L=180.00n
MM2 net9 A2 VDD VNW p18 W=475.00n L=180.00n
MM1 net9 A1 VDD VNW p18 W=475.00n L=180.00n
MM10 ZN B2 net9 VNW p18 W=475.00n L=180.00n
MM0 B2 B2N VDD VNW p18 W=475.00n L=180.00n
MM11 ZN A1 net38 VPW n18 W=280.00n L=180.00n
MM6 ZN B1 net34 VPW n18 W=280.00n L=180.00n
MM12 net34 B2 VSS VPW n18 W=280.00n L=180.00n
MM13 net38 A2 VSS VPW n18 W=280.00n L=180.00n
MM3 B2 B2N VSS VPW n18 W=280.00n L=180.00n
.ENDS AOI22XBUHDV0P4
.SUBCKT AOI22XBUHDV0P7 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM5 ZN B1 net9 VNW p18 W=675.00n L=180.00n
MM2 net9 A2 VDD VNW p18 W=675.00n L=180.00n
MM1 net9 A1 VDD VNW p18 W=675.00n L=180.00n
MM10 ZN B2 net9 VNW p18 W=675.00n L=180.00n
MM0 B2 B2N VDD VNW p18 W=675.00n L=180.00n
MM11 ZN A1 net38 VPW n18 W=560.00n L=180.00n
MM6 ZN B1 net34 VPW n18 W=560.00n L=180.00n
MM12 net34 B2 VSS VPW n18 W=560.00n L=180.00n
MM13 net38 A2 VSS VPW n18 W=560.00n L=180.00n
MM3 B2 B2N VSS VPW n18 W=560.00n L=180.00n
.ENDS AOI22XBUHDV0P7
.SUBCKT AOI22XBUHDV1 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM5 ZN B1 net9 VNW p18 W=1.01u L=180.00n
MM2 net9 A2 VDD VNW p18 W=1.01u L=180.00n
MM1 net9 A1 VDD VNW p18 W=1.01u L=180.00n
MM10 ZN B2 net9 VNW p18 W=1.01u L=180.00n
MM0 B2 B2N VDD VNW p18 W=410.00n L=180.00n
MM11 ZN A1 net38 VPW n18 W=720.00n L=180.00n
MM6 ZN B1 net34 VPW n18 W=720.00n L=180.00n
MM12 net34 B2 VSS VPW n18 W=720.00n L=180.00n
MM13 net38 A2 VSS VPW n18 W=720.00n L=180.00n
MM3 B2 B2N VSS VPW n18 W=290.00n L=180.00n
.ENDS AOI22XBUHDV1
.SUBCKT AOI22XBUHDV2 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM5 ZN B1 net9 VNW p18 W=2.02u L=180.00n
MM2 net9 A2 VDD VNW p18 W=2.02u L=180.00n
MM1 net9 A1 VDD VNW p18 W=2.02u L=180.00n
MM10 ZN B2 net9 VNW p18 W=2.02u L=180.00n
MM0 B2 B2N VDD VNW p18 W=820.00n L=180.00n
MM11 ZN A1 net38 VPW n18 W=1.44u L=180.00n
MM6 ZN B1 net34 VPW n18 W=1.44u L=180.00n
MM12 net34 B2 VSS VPW n18 W=1.44u L=180.00n
MM13 net38 A2 VSS VPW n18 W=1.44u L=180.00n
MM3 B2 B2N VSS VPW n18 W=580.00n L=180.00n
.ENDS AOI22XBUHDV2
.SUBCKT AOI22XBUHDV4 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM5 ZN B1 net9 VNW p18 W=4.04u L=180.00n
MM2 net9 A2 VDD VNW p18 W=3.92u L=180.00n
MM1 net9 A1 VDD VNW p18 W=4.04u L=180.00n
MM10 ZN B2 net9 VNW p18 W=3.93u L=180.00n
MM0 B2 B2N VDD VNW p18 W=1.62u L=180.00n
MM11 ZN A1 net38 VPW n18 W=2.88u L=180.00n
MM6 ZN B1 net34 VPW n18 W=2.88u L=180.00n
MM12 net34 B2 VSS VPW n18 W=2.88u L=180.00n
MM13 net38 A2 VSS VPW n18 W=2.88u L=180.00n
MM3 B2 B2N VSS VPW n18 W=1.16u L=180.00n
.ENDS AOI22XBUHDV4
.SUBCKT AOI2XB11UHDV0P4 A1 A2N B C ZN VDD VSS VNW VPW
MM12 net21 B net026 VNW p18 W=475.000n L=180.00n
MM9 A2 A2N VDD VNW p18 W=475.00n L=180.00n
MM10 net026 A1 VDD VNW p18 W=475.000n L=180.00n
MM11 net026 A2 VDD VNW p18 W=475.000n L=180.00n
MM13 ZN C net21 VNW p18 W=475.000n L=180.00n
MM0 net26 A1 VSS VPW n18 W=280.00n L=180.00n
MM2 ZN B VSS VPW n18 W=280.00n L=180.00n
MM7 ZN C VSS VPW n18 W=280.00n L=180.00n
MM1 ZN A2 net26 VPW n18 W=280.00n L=180.00n
MM8 A2 A2N VSS VPW n18 W=280.00n L=180.00n
.ENDS AOI2XB11UHDV0P4
.SUBCKT AOI2XB11UHDV0P7 A1 A2N B C ZN VDD VSS VNW VPW
MM12 net21 B net026 VNW p18 W=675.000n L=180.00n
MM9 A2 A2N VDD VNW p18 W=410.00n L=180.00n
MM10 net026 A1 VDD VNW p18 W=675.000n L=180.00n
MM11 net026 A2 VDD VNW p18 W=675.000n L=180.00n
MM13 ZN C net21 VNW p18 W=675.000n L=180.00n
MM0 net26 A1 VSS VPW n18 W=560.00n L=180.00n
MM2 ZN B VSS VPW n18 W=560.00n L=180.00n
MM7 ZN C VSS VPW n18 W=560.00n L=180.00n
MM1 ZN A2 net26 VPW n18 W=560.00n L=180.00n
MM8 A2 A2N VSS VPW n18 W=290.00n L=180.00n
.ENDS AOI2XB11UHDV0P7
.SUBCKT AOI2XB11UHDV1 A1 A2N B C ZN VDD VSS VNW VPW
MM12 net21 B net038 VNW p18 W=1.01u L=180.00n
MM9 A2 A2N VDD VNW p18 W=410.00n L=180.00n
MM10 net038 A1 VDD VNW p18 W=1.01u L=180.00n
MM11 net038 A2 VDD VNW p18 W=1.01u L=180.00n
MM13 ZN C net21 VNW p18 W=1.01u L=180.00n
MM0 net26 A1 VSS VPW n18 W=720.00n L=180.00n
MM2 ZN B VSS VPW n18 W=530.00n L=180.00n
MM7 ZN C VSS VPW n18 W=530.00n L=180.00n
MM1 ZN A2 net26 VPW n18 W=720.00n L=180.00n
MM8 A2 A2N VSS VPW n18 W=290.00n L=180.00n
.ENDS AOI2XB11UHDV1
.SUBCKT AOI2XB11UHDV2 A1 A2N B C ZN VDD VSS VNW VPW
MM12 net21 B net038 VNW p18 W=2.02u L=180.00n
MM9 A2 A2N VDD VNW p18 W=820.00n L=180.00n
MM10 net038 A1 VDD VNW p18 W=2.02u L=180.00n
MM11 net038 A2 VDD VNW p18 W=2.02u L=180.00n
MM13 ZN C net21 VNW p18 W=1.95u L=180.00n
MM0 net26 A1 VSS VPW n18 W=1.44u L=180.00n
MM2 ZN B VSS VPW n18 W=1.44u L=180.00n
MM7 ZN C VSS VPW n18 W=1.44u L=180.00n
MM1 ZN A2 net26 VPW n18 W=1.44u L=180.00n
MM8 A2 A2N VSS VPW n18 W=580.00n L=180.00n
.ENDS AOI2XB11UHDV2
.SUBCKT AOI2XB1UHDV0P4 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VDD VNW p18 W=250.00n L=180.00n
MM2 net9 b2n VDD VNW p18 W=400.00n L=180.00n
MM0 net9 B1 VDD VNW p18 W=400.00n L=180.00n
MM1 ZN A net9 VNW p18 W=400.00n L=180.00n
MM6 b2n B2 VSS VPW n18 W=250.00n L=180.00n
MM8 ZN A VSS VPW n18 W=290.00n L=180.00n
MM5 net29 b2n VSS VPW n18 W=290.00n L=180.00n
MM3 ZN B1 net29 VPW n18 W=290.00n L=180.00n
.ENDS AOI2XB1UHDV0P4
.SUBCKT AOI2XB1UHDV0P7 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VDD VNW p18 W=280.00n L=180.00n
MM2 net9 b2n VDD VNW p18 W=710.00n L=180.00n
MM0 net9 B1 VDD VNW p18 W=710.00n L=180.00n
MM1 ZN A net9 VNW p18 W=710.00n L=180.00n
MM6 b2n B2 VSS VPW n18 W=250.00n L=180.00n
MM8 ZN A VSS VPW n18 W=500.00n L=180.00n
MM5 net29 b2n VSS VPW n18 W=500.00n L=180.00n
MM3 ZN B1 net29 VPW n18 W=500.00n L=180.00n
.ENDS AOI2XB1UHDV0P7
.SUBCKT AOI2XB1UHDV1 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VDD VNW p18 W=410.00n L=180.00n
MM2 net9 b2n VDD VNW p18 W=1.01u L=180.00n
MM0 net9 B1 VDD VNW p18 W=1.01u L=180.00n
MM1 ZN A net9 VNW p18 W=1.01u L=180.00n
MM6 b2n B2 VSS VPW n18 W=290.00n L=180.00n
MM8 ZN A VSS VPW n18 W=720.00n L=180.00n
MM5 net29 b2n VSS VPW n18 W=720.00n L=180.00n
MM3 ZN B1 net29 VPW n18 W=720.00n L=180.00n
.ENDS AOI2XB1UHDV1
.SUBCKT AOI2XB1UHDV2 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VDD VNW p18 W=810.00n L=180.00n
MM2 net9 b2n VDD VNW p18 W=2.02u L=180.00n
MM0 net9 B1 VDD VNW p18 W=2.02u L=180.00n
MM1 ZN A net9 VNW p18 W=2.02u L=180.00n
MM6 b2n B2 VSS VPW n18 W=580.00n L=180.00n
MM8 ZN A VSS VPW n18 W=1.44u L=180.00n
MM5 net29 b2n VSS VPW n18 W=1.44u L=180.00n
MM3 ZN B1 net29 VPW n18 W=1.44u L=180.00n
.ENDS AOI2XB1UHDV2
.SUBCKT AOI2XB1UHDV4 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VDD VNW p18 W=1.62u L=180.00n
MM2 net9 b2n VDD VNW p18 W=3.935u L=180.00n
MM0 net9 B1 VDD VNW p18 W=4.04u L=180.00n
MM1 ZN A net9 VNW p18 W=4.04u L=180.00n
MM6 b2n B2 VSS VPW n18 W=1.16u L=180.00n
MM8 ZN A VSS VPW n18 W=2.88u L=180.00n
MM5 net29 b2n VSS VPW n18 W=2.88u L=180.00n
MM3 ZN B1 net29 VPW n18 W=2.88u L=180.00n
.ENDS AOI2XB1UHDV4
.SUBCKT AOI31UHDV0P4 A1 A2 A3 B ZN VDD VSS VNW VPW
MM6 net6 A3 VSS VPW n18 W=0.28u L=180.00n
MM3 ZN A1 net14 VPW n18 W=0.28u L=180.00n
MM5 net14 A2 net6 VPW n18 W=0.28u L=180.00n
MM8 ZN B VSS VPW n18 W=0.28u L=180.00n
MM4 net30 A3 VDD VNW p18 W=490.0n L=180.00n
MM1 ZN B net30 VNW p18 W=490.0n L=180.00n
MM0 net30 A2 VDD VNW p18 W=490.0n L=180.00n
MM2 net30 A1 VDD VNW p18 W=490.0n L=180.00n
.ENDS AOI31UHDV0P4
.SUBCKT AOI31UHDV0P7 A1 A2 A3 B ZN VDD VSS VNW VPW
MM1 ZN B net10 VNW p18 W=0.675u L=180.00n
MM2 net10 A1 VDD VNW p18 W=0.675u L=180.00n
MM0 net10 A2 VDD VNW p18 W=0.675u L=180.00n
MM4 net10 A3 VDD VNW p18 W=0.675u L=180.00n
MM8 ZN B VSS VPW n18 W=560.00n L=180.00n
MM5 net26 A2 net34 VPW n18 W=560.00n L=180.00n
MM3 ZN A1 net26 VPW n18 W=560.00n L=180.00n
MM6 net34 A3 VSS VPW n18 W=560.00n L=180.00n
.ENDS AOI31UHDV0P7
.SUBCKT AOI31UHDV1 A1 A2 A3 B ZN VDD VSS VNW VPW
MM1 ZN B net10 VNW p18 W=1.01u L=180.00n
MM2 net10 A1 VDD VNW p18 W=1.01u L=180.00n
MM0 net10 A2 VDD VNW p18 W=1.01u L=180.00n
MM4 net10 A3 VDD VNW p18 W=1.01u L=180.00n
MM8 ZN B VSS VPW n18 W=720.00n L=180.00n
MM5 net26 A2 net34 VPW n18 W=720.00n L=180.00n
MM3 ZN A1 net26 VPW n18 W=720.00n L=180.00n
MM6 net34 A3 VSS VPW n18 W=720.00n L=180.00n
.ENDS AOI31UHDV1
.SUBCKT AOI31UHDV2 A1 A2 A3 B ZN VDD VSS VNW VPW
MM1 ZN B net10 VNW p18 W=2.02u L=180.00n
MM2 net10 A1 VDD VNW p18 W=2.02u L=180.00n
MM0 net10 A2 VDD VNW p18 W=2.02u L=180.00n
MM4 net10 A3 VDD VNW p18 W=2.02u L=180.00n
MM8 ZN B VSS VPW n18 W=1.44u L=180.00n
MM5 net26 A2 net34 VPW n18 W=1.44u L=180.00n
MM3 ZN A1 net26 VPW n18 W=1000.00n L=180.00n
MM6 net34 A3 VSS VPW n18 W=1.44u L=180.00n
.ENDS AOI31UHDV2
.SUBCKT AOI31UHDV3 A1 A2 A3 B ZN VDD VSS VNW VPW
MM1 ZN B net10 VNW p18 W=3.03u L=180.00n
MM2 net10 A1 VDD VNW p18 W=2.79u L=180.00n
MM0 net10 A2 VDD VNW p18 W=2.87u L=180.00n
MM4 net10 A3 VDD VNW p18 W=3.03u L=180.00n
MM8 ZN B VSS VPW n18 W=2.4u L=180.00n
MM5 net26 A2 net34 VPW n18 W=2.48u L=180.00n
MM3 ZN A1 net26 VPW n18 W=2.56u L=180.00n
MM6 net34 A3 VSS VPW n18 W=2.4u L=180.00n
.ENDS AOI31UHDV3
****Sub-Circuit for AOI32UHDV0P4, Tue Jun  6 11:14:23 CST 2017****
.SUBCKT AOI32UHDV0P4 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM7 net018 B2 VSS VPW n18 W=290.00n L=180.00n
MM8 ZN B1 net018 VPW n18 W=290.00n L=180.00n
MM5 net26 A2 net34 VPW n18 W=290.00n L=180.00n
MM3 ZN A1 net26 VPW n18 W=290.00n L=180.00n
MM6 net34 A3 VSS VPW n18 W=290.00n L=180.00n
MM9 ZN B2 net10 VNW p18 W=490.00n L=180.00n
MM1 ZN B1 net10 VNW p18 W=490.00n L=180.00n
MM2 net10 A1 VDD VNW p18 W=490.00n L=180.00n
MM0 net10 A2 VDD VNW p18 W=490.00n L=180.00n
MM4 net10 A3 VDD VNW p18 W=490.00n L=180.00n
.ENDS AOI32UHDV0P4
****Sub-Circuit for AOI32UHDV0P7, Tue Jun  6 11:14:23 CST 2017****
.SUBCKT AOI32UHDV0P7 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM7 net018 B2 VSS VPW n18 W=560.00n L=180.00n
MM8 ZN B1 net018 VPW n18 W=560.00n L=180.00n
MM5 net26 A2 net34 VPW n18 W=560.00n L=180.00n
MM3 ZN A1 net26 VPW n18 W=560.00n L=180.00n
MM6 net34 A3 VSS VPW n18 W=560.00n L=180.00n
MM9 ZN B2 net10 VNW p18 W=790.00n L=180.00n
MM1 ZN B1 net10 VNW p18 W=790.00n L=180.00n
MM2 net10 A1 VDD VNW p18 W=790.00n L=180.00n
MM0 net10 A2 VDD VNW p18 W=790.00n L=180.00n
MM4 net10 A3 VDD VNW p18 W=790.00n L=180.00n
.ENDS AOI32UHDV0P7
****Sub-Circuit for AOI32UHDV1, Tue Jun  6 11:14:23 CST 2017****
.SUBCKT AOI32UHDV1 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM7 net018 B2 VSS VPW n18 W=720.00n L=180.00n
MM8 ZN B1 net018 VPW n18 W=720.00n L=180.00n
MM5 net26 A2 net34 VPW n18 W=720.00n L=180.00n
MM3 ZN A1 net26 VPW n18 W=720.00n L=180.00n
MM6 net34 A3 VSS VPW n18 W=720.00n L=180.00n
MM9 ZN B2 net10 VNW p18 W=1.01u L=180.00n
MM1 ZN B1 net10 VNW p18 W=1.01u L=180.00n
MM2 net10 A1 VDD VNW p18 W=1.01u L=180.00n
MM0 net10 A2 VDD VNW p18 W=1.01u L=180.00n
MM4 net10 A3 VDD VNW p18 W=1.01u L=180.00n
.ENDS AOI32UHDV1
****Sub-Circuit for AOI32UHDV2, Tue Jun  6 11:14:23 CST 2017****
.SUBCKT AOI32UHDV2 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM7 net018 B2 VSS VPW n18 W=1.44u L=180.00n
MM8 ZN B1 net018 VPW n18 W=1.44u L=180.00n
MM5 net26 A2 net34 VPW n18 W=1.44u L=180.00n
MM3 ZN A1 net26 VPW n18 W=1u L=180.00n
MM6 net34 A3 VSS VPW n18 W=1.44u L=180.00n
MM9 ZN B2 net10 VNW p18 W=2.02u L=180.00n
MM1 ZN B1 net10 VNW p18 W=2.02u L=180.00n
MM2 net10 A1 VDD VNW p18 W=2.02u L=180.00n
MM0 net10 A2 VDD VNW p18 W=2.02u L=180.00n
MM4 net10 A3 VDD VNW p18 W=2.02u L=180.00n
.ENDS AOI32UHDV2
****Sub-Circuit for AOI32UHDV3, Tue Jun  6 11:14:23 CST 2017****
.SUBCKT AOI32UHDV3 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM7 net018 B2 VSS VPW n18 W=2.4u L=180.00n
MM8 ZN B1 net018 VPW n18 W=2.64u L=180.00n
MM5 net26 A2 net34 VPW n18 W=2.48u L=180.00n
MM3 ZN A1 net26 VPW n18 W=2.64u L=180.00n
MM6 net34 A3 VSS VPW n18 W=2.4u L=180.00n
MM9 ZN B2 net10 VNW p18 W=2.95u L=180.00n
MM1 ZN B1 net10 VNW p18 W=2.79u L=180.00n
MM2 net10 A1 VDD VNW p18 W=2.79u L=180.00n
MM0 net10 A2 VDD VNW p18 W=2.87u L=180.00n
MM4 net10 A3 VDD VNW p18 W=3.03u L=180.00n
.ENDS AOI32UHDV3
.SUBCKT BUFUHDV0P4 I Z VDD VSS VNW VPW
MM7 net11 I VDD VNW p18 W=490.00n L=180.00n
MM1 Z net11 VDD VNW p18 W=490.00n L=180.00n
MM15 net11 I VSS VPW n18 W=0.28u L=180.00n
MM0 Z net11 VSS VPW n18 W=0.28u L=180.00n
.ENDS BUFUHDV0P4
.SUBCKT BUFUHDV0P7 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=560.0n L=180.00n
MM15 net7 I VSS VPW n18 W=430.00n L=180.00n
MM1 Z net7 VDD VNW p18 W=790.00n L=180.00n
MM7 net7 I VDD VNW p18 W=500.00n L=180.00n
.ENDS BUFUHDV0P7
.SUBCKT BUFUHDV1 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=720.0n L=180.00n
MM15 net7 I VSS VPW n18 W=430.00n L=180.00n
MM1 Z net7 VDD VNW p18 W=1.01u L=180.00n
MM7 net7 I VDD VNW p18 W=580.00n L=180.00n
.ENDS BUFUHDV1
.SUBCKT BUFUHDV16 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=11.52u L=180.00n
MM15 net7 I VSS VPW n18 W=4.32u L=180.00n
MM1 Z net7 VDD VNW p18 W=16.16u L=180.00n
MM7 net7 I VDD VNW p18 W=6.06u L=180.00n
.ENDS BUFUHDV16
.SUBCKT BUFUHDV2 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=1.44u L=180.00n
MM15 net7 I VSS VPW n18 W=630.00n L=180.00n
MM1 Z net7 VDD VNW p18 W=2.02u L=180.00n
MM7 net7 I VDD VNW p18 W=950.00n L=180.00n
.ENDS BUFUHDV2
.SUBCKT BUFUHDV20 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=14.4u L=180.00n
MM15 net7 I VSS VPW n18 W=5.76u L=180.00n
MM1 Z net7 VDD VNW p18 W=20.2u L=180.00n
MM7 net7 I VDD VNW p18 W=8.08u L=180.00n
.ENDS BUFUHDV20
.SUBCKT BUFUHDV24 I Z VDD VSS VNW VPW
MM7 net11 I VDD VNW p18 W=9.09u L=180.00n
MM1 Z net11 VDD VNW p18 W=24.24u L=180.00n
MM15 net11 I VSS VPW n18 W=6.48u L=180.00n
MM0 Z net11 VSS VPW n18 W=17.28u L=180.00n
.ENDS BUFUHDV24
.SUBCKT BUFUHDV3 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=2.16u L=180.00n
MM15 net7 I VSS VPW n18 W=720.00n L=180.00n
MM1 Z net7 VDD VNW p18 W=3.03u L=180.00n
MM7 net7 I VDD VNW p18 W=1.01u L=180.00n
.ENDS BUFUHDV3
.SUBCKT BUFUHDV4 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=2.88u L=180.00n
MM15 net7 I VSS VPW n18 W=1.12u L=180.00n
MM1 Z net7 VDD VNW p18 W=4.04u L=180.00n
MM7 net7 I VDD VNW p18 W=1.52u L=180.00n
.ENDS BUFUHDV4
.SUBCKT BUFUHDV6 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=4.32u L=180.00n
MM15 net7 I VSS VPW n18 W=1.44u L=180.00n
MM1 Z net7 VDD VNW p18 W=6.06u L=180.00n
MM7 net7 I VDD VNW p18 W=2.02u L=180.00n
.ENDS BUFUHDV6
.SUBCKT BUFUHDV8 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=5.76u L=180.00n
MM15 net7 I VSS VPW n18 W=2.16u L=180.00n
MM1 Z net7 VDD VNW p18 W=8.08u L=180.00n
MM7 net7 I VDD VNW p18 W=3.03u L=180.00n
.ENDS BUFUHDV8
****Sub-Circuit for BUSHOLDUHD, Mon Sep  7 10:31:35 CST 2015****
.SUBCKT BUSHOLDUHD Z VDD VSS VNW VPW
MM2 net031 net10 VDD VNW p18 W=300.00n L=260.00n
MM7 net10 Z VDD VNW p18 W=450.00n L=180.00n
MM1 Z net10 net031 VNW p18 W=300.00n L=260.00n
MM15 net10 Z VSS VPW n18 W=300.00n L=180.00n
MM0 Z net10 net032 VPW n18 W=265.0n L=260.00n
MM3 net032 net10 VSS VPW n18 W=265.0n L=260.00n
.ENDS BUSHOLDUHD
.SUBCKT CLKAND2UHDV0P7 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=0.425u L=180.00n
MM5 net8 A2 VSS VPW n18 W=0.425u L=180.00n
MM3 net24 A1 net8 VPW n18 W=0.425u L=180.00n
MM1 Z net24 VDD VNW p18 W=0.77u L=180.00n
MM0 net24 A2 VDD VNW p18 W=0.475u L=180.00n
MM2 net24 A1 VDD VNW p18 W=0.475u L=180.00n
.ENDS CLKAND2UHDV0P7
.SUBCKT CLKAND2UHDV1 A1 A2 Z VDD VSS VNW VPW
MM2 net4 A1 VDD VNW p18 W=0.465u L=180.00n
MM0 net4 A2 VDD VNW p18 W=0.465u L=180.00n
MM1 Z net4 VDD VNW p18 W=1u L=180.00n
MM3 net4 A1 net20 VPW n18 W=0.425u L=180.00n
MM5 net20 A2 VSS VPW n18 W=0.425u L=180.00n
MM4 Z net4 VSS VPW n18 W=0.425u L=180.00n
.ENDS CLKAND2UHDV1
.SUBCKT CLKAND2UHDV2 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=0.85u L=180.00n
MM5 net8 A2 VSS VPW n18 W=0.425u L=180.00n
MM3 net24 A1 net8 VPW n18 W=0.425u L=180.00n
MM1 Z net24 VDD VNW p18 W=2.02u L=180.00n
MM0 net24 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net24 A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKAND2UHDV2
.SUBCKT CLKAND2UHDV3 A1 A2 Z VDD VSS VNW VPW
MM2 net4 A1 VDD VNW p18 W=1.01u L=180.00n
MM0 net4 A2 VDD VNW p18 W=1.01u L=180.00n
MM1 Z net4 VDD VNW p18 W=3.03u L=180.00n
MM3 net4 A1 net20 VPW n18 W=0.425u L=180.00n
MM5 net20 A2 VSS VPW n18 W=0.425u L=180.00n
MM4 Z net4 VSS VPW n18 W=1.14u L=180.00n
.ENDS CLKAND2UHDV3
.SUBCKT CLKAND2UHDV4 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=1.65u L=180.00n
MM5 net8 A2 VSS VPW n18 W=0.55u L=180.00n
MM3 net24 A1 net8 VPW n18 W=0.55u L=180.00n
MM1 Z net24 VDD VNW p18 W=4.04u L=180.00n
MM0 net24 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net24 A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKAND2UHDV4
.SUBCKT CLKAND2UHDV6 A1 A2 Z VDD VSS VNW VPW
MM4 Z net24 VSS VPW n18 W=2.375u L=180.00n
MM5 net8 A2 VSS VPW n18 W=0.65u L=180.00n
MM3 net24 A1 net8 VPW n18 W=0.65u L=180.00n
MM1 Z net24 VDD VNW p18 W=6.025u L=180.00n
MM0 net24 A2 VDD VNW p18 W=2.02u L=180.00n
MM2 net24 A1 VDD VNW p18 W=2.02u L=180.00n
.ENDS CLKAND2UHDV6
.SUBCKT CLKAND2UHDV8 A1 A2 Z VDD VSS VNW VPW
MM2 net4 A1 VDD VNW p18 W=2.85u L=180.00n
MM0 net4 A2 VDD VNW p18 W=2.97u L=180.00n
MM1 Z net4 VDD VNW p18 W=8.47u L=180.00n
MM3 net4 A1 net20 VPW n18 W=1.17u L=180.00n
MM5 net20 A2 VSS VPW n18 W=1.3u L=180.00n
MM4 Z net4 VSS VPW n18 W=3.12u L=180.00n
.ENDS CLKAND2UHDV8
.SUBCKT CLKBUFUHDV1 I Z VDD VSS VNW VPW
MM15 net3 I VSS VPW n18 W=250.00n L=180.00n
MM0 Z net3 VSS VPW n18 W=320.00n L=180.00n
MM1 Z net3 VDD VNW p18 W=1.01u L=180.00n
MM7 net3 I VDD VNW p18 W=790.00n L=180.00n
.ENDS CLKBUFUHDV1
.SUBCKT CLKBUFUHDV16 I Z VDD VSS VNW VPW
MM15 net11 I VSS VPW n18 W=2.16u L=180.00n
MM0 Z net11 VSS VPW n18 W=5.41u L=180.00n
MM7 net11 I VDD VNW p18 W=6.85u L=180.00n
MM1 Z net11 VDD VNW p18 W=17.13u L=180.00n
.ENDS CLKBUFUHDV16
.SUBCKT CLKBUFUHDV2 I Z VDD VSS VNW VPW
MM0 Z net15 VSS VPW n18 W=600.00n L=180.00n
MM15 net15 I VSS VPW n18 W=250.00n L=180.00n
MM7 net15 I VDD VNW p18 W=840.00n L=180.00n
MM1 Z net15 VDD VNW p18 W=2.02u L=180.00n
.ENDS CLKBUFUHDV2
.SUBCKT CLKBUFUHDV20 I Z VDD VSS VNW VPW
MM15 net11 I VSS VPW n18 W=2.72u L=180.00n
MM0 Z net11 VSS VPW n18 W=6.81u L=180.00n
MM7 net11 I VDD VNW p18 W=8.6u L=180.00n
MM1 Z net11 VDD VNW p18 W=21.49u L=180.00n
.ENDS CLKBUFUHDV20
.SUBCKT CLKBUFUHDV24 I Z VDD VSS VNW VPW
MM0 Z net7 VSS VPW n18 W=7.75u L=180.00n
MM15 net7 I VSS VPW n18 W=3.1u L=180.00n
MM1 Z net7 VDD VNW p18 W=24.46u L=180.00n
MM7 net7 I VDD VNW p18 W=9.78u L=180.00n
.ENDS CLKBUFUHDV24
.SUBCKT CLKBUFUHDV3 I Z VDD VSS VNW VPW
MM15 net3 I VSS VPW n18 W=380.00n L=180.00n
MM0 Z net3 VSS VPW n18 W=1.00u L=180.00n
MM1 Z net3 VDD VNW p18 W=3.03u L=180.00n
MM7 net3 I VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKBUFUHDV3
.SUBCKT CLKBUFUHDV4 I Z VDD VSS VNW VPW
MM15 net7 I VSS VPW n18 W=500.00n L=180.00n
MM0 Z net7 VSS VPW n18 W=1.26u L=180.00n
MM1 Z net7 VDD VNW p18 W=4.04u L=180.00n
MM7 net7 I VDD VNW p18 W=1.62u L=180.00n
.ENDS CLKBUFUHDV4
.SUBCKT CLKBUFUHDV6 I Z VDD VSS VNW VPW
MM0 Z net15 VSS VPW n18 W=1.92u L=180.00n
MM15 net15 I VSS VPW n18 W=700.00n L=180.00n
MM7 net15 I VDD VNW p18 W=2.23u L=180.00n
MM1 Z net15 VDD VNW p18 W=6.06u L=180.00n
.ENDS CLKBUFUHDV6
.SUBCKT CLKBUFUHDV8 I Z VDD VSS VNW VPW
MM15 net11 I VSS VPW n18 W=1.02u L=180.00n
MM0 Z net11 VSS VPW n18 W=2.56u L=180.00n
MM7 net11 I VDD VNW p18 W=3.23u L=180.00n
MM1 Z net11 VDD VNW p18 W=8.08u L=180.00n
.ENDS CLKBUFUHDV8
.SUBCKT CLKINUHDV1 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=320.00n L=180.00n
MM13 ZN I VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKINUHDV1
.SUBCKT CLKINUHDV16 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=5.33u L=180.00n
MM13 ZN I VDD VNW p18 W=16.84u L=180.00n
.ENDS CLKINUHDV16
.SUBCKT CLKINUHDV2 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=600.00n L=180.00n
MM13 ZN I VDD VNW p18 W=2.02u L=180.00n
.ENDS CLKINUHDV2
.SUBCKT CLKINUHDV20 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=6.54u L=180.00n
MM13 ZN I VDD VNW p18 W=20.66u L=180.00n
.ENDS CLKINUHDV20
.SUBCKT CLKINUHDV24 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=7.94u L=180.00n
MM13 ZN I VDD VNW p18 W=25.1u L=180.00n
.ENDS CLKINUHDV24
.SUBCKT CLKINUHDV3 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=1u L=180.00n
MM13 ZN I VDD VNW p18 W=3.03u L=180.00n
.ENDS CLKINUHDV3
.SUBCKT CLKINUHDV4 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=1.26u L=180.00n
MM13 ZN I VDD VNW p18 W=4.04u L=180.00n
.ENDS CLKINUHDV4
.SUBCKT CLKINUHDV6 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=1.9u L=180.00n
MM13 ZN I VDD VNW p18 W=6.01u L=180.00n
.ENDS CLKINUHDV6
.SUBCKT CLKINUHDV8 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=2.66u L=180.00n
MM13 ZN I VDD VNW p18 W=8.41u L=180.00n
.ENDS CLKINUHDV8
.SUBCKT CLKLAHAQUHDV1 CK E Q TE VDD VSS VNW VPW
MM23 ten TE VSS VPW n18 W=420.0n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net77 VSS VPW n18 W=360.0n L=180.00n
MM15 net77 c VSS VPW n18 W=250.00n L=180.00n
MM14 net73 ten VSS VPW n18 W=250.00n L=180.00n
MM13 net77 pm net73 VPW n18 W=250.00n L=180.00n
MM8 pm cn net81 VPW n18 W=0.42u L=180.00n
MM9 net81 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=460.00n L=180.00n
MM5 net93 E VSS VPW n18 W=460.00n L=180.00n
MM4 m pm VSS VPW n18 W=0.42u L=180.00n
MM22 ten TE VDD VNW p18 W=680.0n L=180.00n
MM20 c cn VDD VNW p18 W=520.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net77 VDD VNW p18 W=1.01u L=180.00n
MM12 net28 pm VDD VNW p18 W=810.0n L=180.00n
MM11 net77 c net28 VNW p18 W=810.0n L=180.00n
MM10 net28 ten VDD VNW p18 W=810.0n L=180.00n
MM6 net36 m VDD VNW p18 W=415.000n L=180.00n
MM7 pm c net36 VNW p18 W=415.000n L=180.00n
MM2 net48 E VDD VNW p18 W=680.0n L=180.00n
MM0 pm cn net48 VNW p18 W=680.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHAQUHDV1
.SUBCKT CLKLAHAQUHDV2 CK E Q TE VDD VSS VNW VPW
MM4 m pm VSS VPW n18 W=400.0n L=180.00n
MM5 net9 E VSS VPW n18 W=540.00n L=180.00n
MM3 pm c net9 VPW n18 W=540.00n L=180.00n
MM9 net17 m VSS VPW n18 W=0.42u L=180.00n
MM8 pm cn net17 VPW n18 W=0.42u L=180.00n
MM13 net25 pm net29 VPW n18 W=430.00n L=180.00n
MM14 net29 ten VSS VPW n18 W=430.00n L=180.00n
MM15 net25 c VSS VPW n18 W=430.00n L=180.00n
MM17 Q net25 VSS VPW n18 W=740.00n L=180.00n
MM19 cn CK VSS VPW n18 W=570.0n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM23 ten TE VSS VPW n18 W=460.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
MM0 pm cn net60 VNW p18 W=810.0n L=180.00n
MM2 net60 E VDD VNW p18 W=810.0n L=180.00n
MM7 pm c net68 VNW p18 W=0.415u L=180.00n
MM6 net68 m VDD VNW p18 W=0.415u L=180.00n
MM10 net80 ten VDD VNW p18 W=1.82u L=180.00n
MM11 net25 c net80 VNW p18 W=1.82u L=180.00n
MM12 net80 pm VDD VNW p18 W=1.82u L=180.00n
MM16 Q net25 VDD VNW p18 W=2.02u L=180.00n
MM18 cn CK VDD VNW p18 W=870.0n L=180.00n
MM20 c cn VDD VNW p18 W=870.0n L=180.00n
MM22 ten TE VDD VNW p18 W=680.0n L=180.00n
.ENDS CLKLAHAQUHDV2
.SUBCKT CLKLAHAQUHDV3 CK E Q TE VDD VSS VNW VPW
MM4 m pm VSS VPW n18 W=400.0n L=180.00n
MM5 net9 E VSS VPW n18 W=540.00n L=180.00n
MM3 pm c net9 VPW n18 W=540.00n L=180.00n
MM9 net17 m VSS VPW n18 W=0.42u L=180.00n
MM8 pm cn net17 VPW n18 W=0.42u L=180.00n
MM13 net25 pm net29 VPW n18 W=430.00n L=180.00n
MM14 net29 ten VSS VPW n18 W=430.00n L=180.00n
MM15 net25 c VSS VPW n18 W=430.00n L=180.00n
MM17 Q net25 VSS VPW n18 W=1.15u L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM21 c cn VSS VPW n18 W=420.0n L=180.00n
MM23 ten TE VSS VPW n18 W=460.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
MM0 pm cn net60 VNW p18 W=0.85u L=180.00n
MM2 net60 E VDD VNW p18 W=810.0n L=180.00n
MM7 pm c net68 VNW p18 W=0.415u L=180.00n
MM6 net68 m VDD VNW p18 W=0.415u L=180.00n
MM10 net80 ten VDD VNW p18 W=1.82u L=180.00n
MM11 net25 c net80 VNW p18 W=1.82u L=180.00n
MM12 net80 pm VDD VNW p18 W=1.82u L=180.00n
MM16 Q net25 VDD VNW p18 W=3.03u L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM20 c cn VDD VNW p18 W=680.0n L=180.00n
MM22 ten TE VDD VNW p18 W=680.0n L=180.00n
.ENDS CLKLAHAQUHDV3
.SUBCKT CLKLAHAQUHDV4 CK E Q TE VDD VSS VNW VPW
MM23 ten TE VSS VPW n18 W=430.0n L=180.00n
MM21 c cn VSS VPW n18 W=420.0n L=180.00n
MM19 cn CK VSS VPW n18 W=570.0n L=180.00n
MM17 Q net77 VSS VPW n18 W=1.56u L=180.00n
MM15 net77 c VSS VPW n18 W=430.00n L=180.00n
MM14 net73 ten VSS VPW n18 W=430.00n L=180.00n
MM13 net77 pm net73 VPW n18 W=430.00n L=180.00n
MM8 pm cn net85 VPW n18 W=0.42u L=180.00n
MM9 net85 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=570.00n L=180.00n
MM5 net93 E VSS VPW n18 W=570.00n L=180.00n
MM4 m pm VSS VPW n18 W=400.0n L=180.00n
MM22 ten TE VDD VNW p18 W=680.0n L=180.00n
MM20 c cn VDD VNW p18 W=870.0n L=180.00n
MM18 cn CK VDD VNW p18 W=870.0n L=180.00n
MM16 Q net77 VDD VNW p18 W=4.04u L=180.00n
MM12 net28 pm VDD VNW p18 W=1.82u L=180.00n
MM11 net77 c net28 VNW p18 W=1.82u L=180.00n
MM10 net28 ten VDD VNW p18 W=1.82u L=180.00n
MM6 net40 m VDD VNW p18 W=0.415u L=180.00n
MM7 pm c net40 VNW p18 W=0.415u L=180.00n
MM2 net48 E VDD VNW p18 W=0.81u L=180.00n
MM0 pm cn net48 VNW p18 W=850.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHAQUHDV4
.SUBCKT CLKLAHAQUHDV6 CK E Q TE VDD VSS VNW VPW
MM23 ten TE VSS VPW n18 W=0.545u L=180.00n
MM21 c cn VSS VPW n18 W=420.0n L=180.00n
MM19 cn CK VSS VPW n18 W=570.0n L=180.00n
MM17 Q net77 VSS VPW n18 W=2.29u L=180.00n
MM15 net77 c VSS VPW n18 W=860.0n L=180.00n
MM14 net73 ten VSS VPW n18 W=860.0n L=180.00n
MM13 net77 pm net73 VPW n18 W=860.0n L=180.00n
MM8 pm cn net85 VPW n18 W=0.42u L=180.00n
MM9 net85 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=570.00n L=180.00n
MM5 net93 E VSS VPW n18 W=570.00n L=180.00n
MM4 m pm VSS VPW n18 W=400.0n L=180.00n
MM22 ten TE VDD VNW p18 W=0.835u L=180.00n
MM20 c cn VDD VNW p18 W=870.0n L=180.00n
MM18 cn CK VDD VNW p18 W=870.0n L=180.00n
MM16 Q net77 VDD VNW p18 W=6.06u L=180.00n
MM12 net28 pm VDD VNW p18 W=3.64u L=180.00n
MM11 net77 c net28 VNW p18 W=3.64u L=180.00n
MM10 net28 ten VDD VNW p18 W=3.64u L=180.00n
MM6 net40 m VDD VNW p18 W=0.415u L=180.00n
MM7 pm c net40 VNW p18 W=0.415u L=180.00n
MM2 net48 E VDD VNW p18 W=0.81u L=180.00n
MM0 pm cn net48 VNW p18 W=850.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHAQUHDV6
.SUBCKT CLKLAHAQUHDV8 CK E Q TE VDD VSS VNW VPW
MM23 ten TE VSS VPW n18 W=0.545u L=180.00n
MM21 c cn VSS VPW n18 W=420.0n L=180.00n
MM19 cn CK VSS VPW n18 W=570.0n L=180.00n
MM17 Q net77 VSS VPW n18 W=3.09u L=180.00n
MM15 net77 c VSS VPW n18 W=860.0n L=180.00n
MM14 net73 ten VSS VPW n18 W=860.0n L=180.00n
MM13 net77 pm net73 VPW n18 W=860.0n L=180.00n
MM8 pm cn net85 VPW n18 W=0.42u L=180.00n
MM9 net85 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=570.00n L=180.00n
MM5 net93 E VSS VPW n18 W=570.00n L=180.00n
MM4 m pm VSS VPW n18 W=400.0n L=180.00n
MM22 ten TE VDD VNW p18 W=0.835u L=180.00n
MM20 c cn VDD VNW p18 W=870.0n L=180.00n
MM18 cn CK VDD VNW p18 W=870.0n L=180.00n
MM16 Q net77 VDD VNW p18 W=8.08u L=180.00n
MM12 net28 pm VDD VNW p18 W=3.64u L=180.00n
MM11 net77 c net28 VNW p18 W=3.64u L=180.00n
MM10 net28 ten VDD VNW p18 W=3.64u L=180.00n
MM6 net40 m VDD VNW p18 W=0.415u L=180.00n
MM7 pm c net40 VNW p18 W=0.415u L=180.00n
MM2 net48 E VDD VNW p18 W=0.81u L=180.00n
MM0 pm cn net48 VNW p18 W=850.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHAQUHDV8
****Sub-Circuit for CLKLAHQUHDV1, Tue Jun 13 16:51:01 CST 2017****
.SUBCKT CLKLAHQUHDV1 CK E Q TE VDD VSS VNW VPW
MM14 net93 TE VSS VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net77 VSS VPW n18 W=320.0n L=180.00n
MM15 net77 c VSS VPW n18 W=250.00n L=180.00n
MM13 net77 pm VSS VPW n18 W=250.00n L=180.00n
MM8 pm cn net81 VPW n18 W=0.42u L=180.00n
MM9 net81 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=460.00n L=180.00n
MM5 net93 E VSS VPW n18 W=460.00n L=180.00n
MM4 m pm VSS VPW n18 W=0.42u L=180.00n
MM20 c cn VDD VNW p18 W=520.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net77 VDD VNW p18 W=1.01u L=180.00n
MM12 net28 pm VDD VNW p18 W=410.0n L=180.00n
MM11 net77 c net28 VNW p18 W=410.0n L=180.00n
MM6 net36 m VDD VNW p18 W=415.000n L=180.00n
MM7 pm c net36 VNW p18 W=415.000n L=180.00n
MM2 net48 E net0159 VNW p18 W=680.0n L=180.00n
MM10 net0159 TE VDD VNW p18 W=680.0n L=180.00n
MM0 pm cn net48 VNW p18 W=680.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHQUHDV1
****Sub-Circuit for CLKLAHQUHDV2, Tue Jun 13 16:51:01 CST 2017****
.SUBCKT CLKLAHQUHDV2 CK E Q TE VDD VSS VNW VPW
MM14 net93 TE VSS VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q pq VSS VPW n18 W=830.0n L=180.00n
MM15 pq c VSS VPW n18 W=250.00n L=180.00n
MM13 pq pm VSS VPW n18 W=250.00n L=180.00n
MM8 pm cn net81 VPW n18 W=0.42u L=180.00n
MM9 net81 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=460.00n L=180.00n
MM5 net93 E VSS VPW n18 W=460.00n L=180.00n
MM4 m pm VSS VPW n18 W=0.42u L=180.00n
MM20 c cn VDD VNW p18 W=520.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q pq VDD VNW p18 W=2.02u L=180.00n
MM12 net28 pm VDD VNW p18 W=1.01u L=180.00n
MM11 pq c net28 VNW p18 W=1.01u L=180.00n
MM6 net36 m VDD VNW p18 W=415.000n L=180.00n
MM7 pm c net36 VNW p18 W=415.000n L=180.00n
MM2 net48 E net0159 VNW p18 W=680.0n L=180.00n
MM10 net0159 TE VDD VNW p18 W=680.0n L=180.00n
MM0 pm cn net48 VNW p18 W=680.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHQUHDV2
****Sub-Circuit for CLKLAHQUHDV3, Tue Jun 13 16:51:01 CST 2017****
.SUBCKT CLKLAHQUHDV3 CK E Q TE VDD VSS VNW VPW
MM14 net93 TE VSS VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q pq VSS VPW n18 W=1.3u L=180.00n
MM15 pq c VSS VPW n18 W=250.00n L=180.00n
MM13 pq pm VSS VPW n18 W=250.00n L=180.00n
MM8 pm cn net81 VPW n18 W=0.42u L=180.00n
MM9 net81 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=460.00n L=180.00n
MM5 net93 E VSS VPW n18 W=460.00n L=180.00n
MM4 m pm VSS VPW n18 W=0.42u L=180.00n
MM20 c cn VDD VNW p18 W=520.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q pq VDD VNW p18 W=3.03u L=180.00n
MM12 net28 pm VDD VNW p18 W=1.01u L=180.00n
MM11 pq c net28 VNW p18 W=1.01u L=180.00n
MM6 net36 m VDD VNW p18 W=415.000n L=180.00n
MM7 pm c net36 VNW p18 W=415.000n L=180.00n
MM2 net48 E net0159 VNW p18 W=680.0n L=180.00n
MM10 net0159 TE VDD VNW p18 W=680.0n L=180.00n
MM0 pm cn net48 VNW p18 W=680.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHQUHDV3
****Sub-Circuit for CLKLAHQUHDV4, Tue Jun 13 16:51:01 CST 2017****
.SUBCKT CLKLAHQUHDV4 CK E Q TE VDD VSS VNW VPW
MM14 net93 TE VSS VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q pq VSS VPW n18 W=1.77u L=180.00n
MM15 pq c VSS VPW n18 W=400.00n L=180.00n
MM13 pq pm VSS VPW n18 W=400.00n L=180.00n
MM8 pm cn net81 VPW n18 W=0.42u L=180.00n
MM9 net81 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=460.00n L=180.00n
MM5 net93 E VSS VPW n18 W=460.00n L=180.00n
MM4 m pm VSS VPW n18 W=0.42u L=180.00n
MM20 c cn VDD VNW p18 W=520.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q pq VDD VNW p18 W=4.04u L=180.00n
MM12 net28 pm VDD VNW p18 W=1.61u L=180.00n
MM11 pq c net28 VNW p18 W=1.61u L=180.00n
MM6 net36 m VDD VNW p18 W=415.000n L=180.00n
MM7 pm c net36 VNW p18 W=415.000n L=180.00n
MM2 net48 E net0159 VNW p18 W=680.0n L=180.00n
MM10 net0159 TE VDD VNW p18 W=680.0n L=180.00n
MM0 pm cn net48 VNW p18 W=680.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHQUHDV4
****Sub-Circuit for CLKLAHQUHDV6, Tue Jun 13 16:59:42 CST 2017****
.SUBCKT CLKLAHQUHDV6 CK E Q TE VDD VSS VNW VPW
MM14 net93 TE VSS VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q pq VSS VPW n18 W=2.59u L=180.00n
MM15 pq c VSS VPW n18 W=420.00n L=180.00n
MM13 pq pm VSS VPW n18 W=420.00n L=180.00n
MM8 pm cn net81 VPW n18 W=0.42u L=180.00n
MM9 net81 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=460.00n L=180.00n
MM5 net93 E VSS VPW n18 W=460.00n L=180.00n
MM4 m pm VSS VPW n18 W=0.42u L=180.00n
MM20 c cn VDD VNW p18 W=520.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q pq VDD VNW p18 W=6.06u L=180.00n
MM12 net28 pm VDD VNW p18 W=2.02u L=180.00n
MM11 pq c net28 VNW p18 W=2.02u L=180.00n
MM6 net36 m VDD VNW p18 W=415.000n L=180.00n
MM7 pm c net36 VNW p18 W=415.000n L=180.00n
MM2 net48 E net0159 VNW p18 W=680.0n L=180.00n
MM10 net0159 TE VDD VNW p18 W=680.0n L=180.00n
MM0 pm cn net48 VNW p18 W=680.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHQUHDV6
****Sub-Circuit for CLKLAHQUHDV8, Tue Jun 13 16:51:01 CST 2017****
.SUBCKT CLKLAHQUHDV8 CK E Q TE VDD VSS VNW VPW
MM14 net93 TE VSS VPW n18 W=570.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q pq VSS VPW n18 W=3.41u L=180.00n
MM15 pq c VSS VPW n18 W=800.0n L=180.00n
MM13 pq pm VSS VPW n18 W=800.0n L=180.00n
MM8 pm cn net81 VPW n18 W=0.42u L=180.00n
MM9 net81 m VSS VPW n18 W=0.42u L=180.00n
MM3 pm c net93 VPW n18 W=570.00n L=180.00n
MM5 net93 E VSS VPW n18 W=570.00n L=180.00n
MM4 m pm VSS VPW n18 W=0.42u L=180.00n
MM20 c cn VDD VNW p18 W=520.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q pq VDD VNW p18 W=8.08u L=180.00n
MM12 net28 pm VDD VNW p18 W=2.965u L=180.00n
MM11 pq c net28 VNW p18 W=2.965u L=180.00n
MM6 net36 m VDD VNW p18 W=415.000n L=180.00n
MM7 pm c net36 VNW p18 W=415.000n L=180.00n
MM2 net48 E net0159 VNW p18 W=810.0n L=180.00n
MM10 net0159 TE VDD VNW p18 W=810.0n L=180.00n
MM0 pm cn net48 VNW p18 W=810.0n L=180.00n
MM1 m pm VDD VNW p18 W=0.42u L=180.00n
.ENDS CLKLAHQUHDV8
****Sub-Circuit for CLKLANAQUHDV1, Tue Jun 13 17:49:43 CST 2017****
.SUBCKT CLKLANAQUHDV1 CK E Q TE VDD VSS VNW VPW
MM25 net0215 E VSS VPW n18 W=460.00n L=180.00n
MM3 pm cn net0215 VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net69 VSS VPW n18 W=420.0n L=180.00n
MM14 net65 m VSS VPW n18 W=540.00n L=180.00n
MM13 net69 c net65 VPW n18 W=720.00n L=180.00n
MM8 pm c net77 VPW n18 W=0.43u L=180.00n
MM9 net77 m VSS VPW n18 W=0.43u L=180.00n
MM22 net65 TE VSS VPW n18 W=720.00n L=180.00n
MM4 m pm VSS VPW n18 W=460.0n L=180.00n
MM0 pm c net0174 VNW p18 W=810.0n L=180.00n
MM2 net0174 E VDD VNW p18 W=810.0n L=180.00n
MM15 net0149 TE VDD VNW p18 W=0.42u L=180.00n
MM20 c cn VDD VNW p18 W=420.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net69 VDD VNW p18 W=1.01u L=180.00n
MM12 net69 c VDD VNW p18 W=0.42u L=180.00n
MM11 net69 m net0149 VNW p18 W=0.42u L=180.00n
MM6 net36 m VDD VNW p18 W=0.44u L=180.00n
MM7 pm cn net36 VNW p18 W=0.44u L=180.00n
MM1 m pm VDD VNW p18 W=580.00n L=180.00n
.ENDS CLKLANAQUHDV1
****Sub-Circuit for CLKLANAQUHDV2, Tue Jun 13 17:49:43 CST 2017****
.SUBCKT CLKLANAQUHDV2 CK E Q TE VDD VSS VNW VPW
MM25 net0215 E VSS VPW n18 W=460.00n L=180.00n
MM3 pm cn net0215 VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net69 VSS VPW n18 W=720.0n L=180.00n
MM14 net65 m VSS VPW n18 W=540.00n L=180.00n
MM13 net69 c net65 VPW n18 W=540.00n L=180.00n
MM8 pm c net77 VPW n18 W=0.43u L=180.00n
MM9 net77 m VSS VPW n18 W=0.43u L=180.00n
MM22 net65 TE VSS VPW n18 W=540.00n L=180.00n
MM4 m pm VSS VPW n18 W=460.0n L=180.00n
MM0 pm c net0174 VNW p18 W=810.0n L=180.00n
MM2 net0174 E VDD VNW p18 W=810.0n L=180.00n
MM15 net0149 TE VDD VNW p18 W=810.00n L=180.00n
MM20 c cn VDD VNW p18 W=420.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net69 VDD VNW p18 W=2.02u L=180.00n
MM12 net69 c VDD VNW p18 W=810.00n L=180.00n
MM11 net69 m net0149 VNW p18 W=810.00n L=180.00n
MM6 net36 m VDD VNW p18 W=0.44u L=180.00n
MM7 pm cn net36 VNW p18 W=0.44u L=180.00n
MM1 m pm VDD VNW p18 W=580.00n L=180.00n
.ENDS CLKLANAQUHDV2
****Sub-Circuit for CLKLANAQUHDV3, Tue Jun 13 17:49:43 CST 2017****
.SUBCKT CLKLANAQUHDV3 CK E Q TE VDD VSS VNW VPW
MM25 net0215 E VSS VPW n18 W=460.00n L=180.00n
MM3 pm cn net0215 VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net69 VSS VPW n18 W=1.08u L=180.00n
MM14 net65 m VSS VPW n18 W=540.00n L=180.00n
MM13 net69 c net65 VPW n18 W=700.00n L=180.00n
MM8 pm c net77 VPW n18 W=0.43u L=180.00n
MM9 net77 m VSS VPW n18 W=0.43u L=180.00n
MM22 net65 TE VSS VPW n18 W=700.00n L=180.00n
MM4 m pm VSS VPW n18 W=460.0n L=180.00n
MM0 pm c net0174 VNW p18 W=810.0n L=180.00n
MM2 net0174 E VDD VNW p18 W=810.0n L=180.00n
MM15 net0149 TE VDD VNW p18 W=920.00n L=180.00n
MM20 c cn VDD VNW p18 W=420.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net69 VDD VNW p18 W=3.03u L=180.00n
MM12 net69 c VDD VNW p18 W=920.00n L=180.00n
MM11 net69 m net0149 VNW p18 W=920.00n L=180.00n
MM6 net36 m VDD VNW p18 W=0.44u L=180.00n
MM7 pm cn net36 VNW p18 W=0.44u L=180.00n
MM1 m pm VDD VNW p18 W=580.00n L=180.00n
.ENDS CLKLANAQUHDV3
****Sub-Circuit for CLKLANAQUHDV4, Tue Jun 13 17:49:43 CST 2017****
.SUBCKT CLKLANAQUHDV4 CK E Q TE VDD VSS VNW VPW
MM25 net0215 E VSS VPW n18 W=460.00n L=180.00n
MM3 pm cn net0215 VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net69 VSS VPW n18 W=1.44u L=180.00n
MM14 net65 m VSS VPW n18 W=1.08u L=180.00n
MM13 net69 c net65 VPW n18 W=1.08u L=180.00n
MM8 pm c net77 VPW n18 W=0.43u L=180.00n
MM9 net77 m VSS VPW n18 W=0.43u L=180.00n
MM22 net65 TE VSS VPW n18 W=1.08u L=180.00n
MM4 m pm VSS VPW n18 W=460.0n L=180.00n
MM0 pm c net0174 VNW p18 W=810.0n L=180.00n
MM2 net0174 E VDD VNW p18 W=810.0n L=180.00n
MM15 net0149 TE VDD VNW p18 W=1.62u L=180.00n
MM20 c cn VDD VNW p18 W=420.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net69 VDD VNW p18 W=4.04u L=180.00n
MM12 net69 c VDD VNW p18 W=1.62u L=180.00n
MM11 net69 m net0149 VNW p18 W=1.62u L=180.00n
MM6 net36 m VDD VNW p18 W=0.44u L=180.00n
MM7 pm cn net36 VNW p18 W=0.44u L=180.00n
MM1 m pm VDD VNW p18 W=580.00n L=180.00n
.ENDS CLKLANAQUHDV4
****Sub-Circuit for CLKLANAQUHDV6, Tue Jun 13 17:49:43 CST 2017****
.SUBCKT CLKLANAQUHDV6 CK E Q TE VDD VSS VNW VPW
MM25 net0215 E VSS VPW n18 W=460.00n L=180.00n
MM3 pm cn net0215 VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net69 VSS VPW n18 W=2.16u L=180.00n
MM14 net65 m VSS VPW n18 W=1.08u L=180.00n
MM13 net69 c net65 VPW n18 W=1.14u L=180.00n
MM8 pm c net77 VPW n18 W=0.43u L=180.00n
MM9 net77 m VSS VPW n18 W=0.43u L=180.00n
MM22 net65 TE VSS VPW n18 W=1.08u L=180.00n
MM4 m pm VSS VPW n18 W=560.0n L=180.00n
MM0 pm c net0174 VNW p18 W=810.0n L=180.00n
MM2 net0174 E VDD VNW p18 W=810.0n L=180.00n
MM15 net0149 TE VDD VNW p18 W=1.84u L=180.00n
MM20 c cn VDD VNW p18 W=420.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net69 VDD VNW p18 W=6.05u L=180.00n
MM12 net69 c VDD VNW p18 W=2.42u L=180.00n
MM11 net69 m net0149 VNW p18 W=1.84u L=180.00n
MM6 net36 m VDD VNW p18 W=0.44u L=180.00n
MM7 pm cn net36 VNW p18 W=0.44u L=180.00n
MM1 m pm VDD VNW p18 W=730.00n L=180.00n
.ENDS CLKLANAQUHDV6
****Sub-Circuit for CLKLANAQUHDV8, Tue Jun 13 17:49:43 CST 2017****
.SUBCKT CLKLANAQUHDV8 CK E Q TE VDD VSS VNW VPW
MM25 net0215 E VSS VPW n18 W=460.00n L=180.00n
MM3 pm cn net0215 VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net69 VSS VPW n18 W=2.88u L=180.00n
MM14 net65 m VSS VPW n18 W=1.7u L=180.00n
MM13 net69 c net65 VPW n18 W=1.7u L=180.00n
MM8 pm c net77 VPW n18 W=0.43u L=180.00n
MM9 net77 m VSS VPW n18 W=0.43u L=180.00n
MM22 net65 TE VSS VPW n18 W=1.62u L=180.00n
MM4 m pm VSS VPW n18 W=670.00n L=180.00n
MM0 pm c net0174 VNW p18 W=810.0n L=180.00n
MM2 net0174 E VDD VNW p18 W=810.0n L=180.00n
MM15 net0149 TE VDD VNW p18 W=1.84u L=180.00n
MM20 c cn VDD VNW p18 W=420.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net69 VDD VNW p18 W=7.57u L=180.00n
MM12 net69 c VDD VNW p18 W=3.24u L=180.00n
MM11 net69 m net0149 VNW p18 W=1.84u L=180.00n
MM6 net36 m VDD VNW p18 W=0.44u L=180.00n
MM7 pm cn net36 VNW p18 W=0.44u L=180.00n
MM1 m pm VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKLANAQUHDV8
.SUBCKT CLKLANQUHDV1 CK E Q TE VDD VSS VNW VPW
MM25 net0215 E VSS VPW n18 W=460.00n L=180.00n
MM3 pm cn net0215 VPW n18 W=460.00n L=180.00n
MM5 net0215 TE VSS VPW n18 W=460.00n L=180.00n
MM21 c cn VSS VPW n18 W=460.0n L=180.00n
MM19 cn CK VSS VPW n18 W=460.0n L=180.00n
MM17 Q net69 VSS VPW n18 W=410.0n L=180.00n
MM14 net65 m VSS VPW n18 W=720.00n L=180.00n
MM13 net69 c net65 VPW n18 W=720.00n L=180.00n
MM8 pm c net77 VPW n18 W=0.43u L=180.00n
MM9 net77 m VSS VPW n18 W=0.43u L=180.00n
MM4 m pm VSS VPW n18 W=460.0n L=180.00n
MM24 net0170 TE VDD VNW p18 W=810.0n L=180.00n
MM0 pm c net0174 VNW p18 W=810.0n L=180.00n
MM2 net0174 E net0170 VNW p18 W=810.0n L=180.00n
MM20 c cn VDD VNW p18 W=420.0n L=180.00n
MM18 cn CK VDD VNW p18 W=680.0n L=180.00n
MM16 Q net69 VDD VNW p18 W=1.01u L=180.00n
MM12 net69 c VDD VNW p18 W=0.42u L=180.00n
MM11 net69 m VDD VNW p18 W=0.42u L=180.00n
MM6 net36 m VDD VNW p18 W=0.44u L=180.00n
MM7 pm cn net36 VNW p18 W=0.44u L=180.00n
MM1 m pm VDD VNW p18 W=580.00n L=180.00n
.ENDS CLKLANQUHDV1
.SUBCKT CLKLANQUHDV2 CK E Q TE VDD VSS VNW VPW
MM4 m pm VSS VPW n18 W=0.47u L=180.00n
MM9 net9 m VSS VPW n18 W=0.43u L=180.00n
MM8 pm c net9 VPW n18 W=0.43u L=180.00n
MM13 net17 c net21 VPW n18 W=720.00n L=180.00n
MM14 net21 m VSS VPW n18 W=720.00n L=180.00n
MM17 Q net17 VSS VPW n18 W=730.00n L=180.00n
MM25 net33 E VSS VPW n18 W=0.47u L=180.00n
MM5 net33 TE VSS VPW n18 W=0.47u L=180.00n
MM3 pm cn net33 VPW n18 W=0.47u L=180.00n
MM19 cn CK VSS VPW n18 W=0.58u L=180.00n
MM21 c cn VSS VPW n18 W=0.58u L=180.00n
MM1 m pm VDD VNW p18 W=0.69u L=180.00n
MM7 pm cn net56 VNW p18 W=0.42u L=180.00n
MM6 net56 m VDD VNW p18 W=0.42u L=180.00n
MM11 net17 m VDD VNW p18 W=1.01u L=180.00n
MM12 net17 c VDD VNW p18 W=1.01u L=180.00n
MM16 Q net17 VDD VNW p18 W=2.02u L=180.00n
MM24 net84 TE VDD VNW p18 W=0.975u L=180.00n
MM0 pm c net80 VNW p18 W=0.975u L=180.00n
MM2 net80 E net84 VNW p18 W=0.975u L=180.00n
MM18 cn CK VDD VNW p18 W=0.88u L=180.00n
MM20 c cn VDD VNW p18 W=750.00n L=180.00n
.ENDS CLKLANQUHDV2
.SUBCKT CLKLANQUHDV3 CK E Q TE VDD VSS VNW VPW
MM4 m pm VSS VPW n18 W=0.47u L=180.00n
MM9 net9 m VSS VPW n18 W=0.43u L=180.00n
MM8 pm c net9 VPW n18 W=0.43u L=180.00n
MM13 net17 c net21 VPW n18 W=720.00n L=180.00n
MM14 net21 m VSS VPW n18 W=720.00n L=180.00n
MM17 Q net17 VSS VPW n18 W=1.14u L=180.00n
MM25 net33 E VSS VPW n18 W=0.47u L=180.00n
MM5 net33 TE VSS VPW n18 W=0.47u L=180.00n
MM3 pm cn net33 VPW n18 W=0.47u L=180.00n
MM19 cn CK VSS VPW n18 W=0.58u L=180.00n
MM21 c cn VSS VPW n18 W=0.58u L=180.00n
MM1 m pm VDD VNW p18 W=0.69u L=180.00n
MM7 pm cn net56 VNW p18 W=0.42u L=180.00n
MM6 net56 m VDD VNW p18 W=0.42u L=180.00n
MM11 net17 m VDD VNW p18 W=1.01u L=180.00n
MM12 net17 c VDD VNW p18 W=1.01u L=180.00n
MM16 Q net17 VDD VNW p18 W=3.03u L=180.00n
MM24 net84 TE VDD VNW p18 W=0.975u L=180.00n
MM0 pm c net80 VNW p18 W=0.975u L=180.00n
MM2 net80 E net84 VNW p18 W=0.975u L=180.00n
MM18 cn CK VDD VNW p18 W=0.88u L=180.00n
MM20 c cn VDD VNW p18 W=750.00n L=180.00n
.ENDS CLKLANQUHDV3
.SUBCKT CLKLANQUHDV4 CK E Q TE VDD VSS VNW VPW
MM4 m pm VSS VPW n18 W=0.47u L=180.00n
MM9 net9 m VSS VPW n18 W=0.43u L=180.00n
MM8 pm c net9 VPW n18 W=0.43u L=180.00n
MM13 net17 c net21 VPW n18 W=720.00n L=180.00n
MM14 net21 m VSS VPW n18 W=720.00n L=180.00n
MM17 Q net17 VSS VPW n18 W=1.55u L=180.00n
MM25 net33 E VSS VPW n18 W=0.47u L=180.00n
MM5 net33 TE VSS VPW n18 W=0.47u L=180.00n
MM3 pm cn net33 VPW n18 W=0.47u L=180.00n
MM19 cn CK VSS VPW n18 W=0.58u L=180.00n
MM21 c cn VSS VPW n18 W=0.58u L=180.00n
MM1 m pm VDD VNW p18 W=0.69u L=180.00n
MM7 pm cn net56 VNW p18 W=0.42u L=180.00n
MM6 net56 m VDD VNW p18 W=0.42u L=180.00n
MM11 net17 m VDD VNW p18 W=1.01u L=180.00n
MM12 net17 c VDD VNW p18 W=1.01u L=180.00n
MM16 Q net17 VDD VNW p18 W=4.04u L=180.00n
MM24 net84 TE VDD VNW p18 W=0.975u L=180.00n
MM0 pm c net80 VNW p18 W=0.975u L=180.00n
MM2 net80 E net84 VNW p18 W=0.975u L=180.00n
MM18 cn CK VDD VNW p18 W=0.88u L=180.00n
MM20 c cn VDD VNW p18 W=750.00n L=180.00n
.ENDS CLKLANQUHDV4
.SUBCKT CLKLANQUHDV6 CK E Q TE VDD VSS VNW VPW
MM4 m pm VSS VPW n18 W=0.47u L=180.00n
MM9 net9 m VSS VPW n18 W=0.43u L=180.00n
MM8 pm c net9 VPW n18 W=0.43u L=180.00n
MM13 net17 c net21 VPW n18 W=1.44u L=180.00n
MM14 net21 m VSS VPW n18 W=1.44u L=180.00n
MM17 Q net17 VSS VPW n18 W=2.3u L=180.00n
MM25 net33 E VSS VPW n18 W=0.47u L=180.00n
MM5 net33 TE VSS VPW n18 W=0.47u L=180.00n
MM3 pm cn net33 VPW n18 W=0.47u L=180.00n
MM19 cn CK VSS VPW n18 W=0.58u L=180.00n
MM21 c cn VSS VPW n18 W=0.58u L=180.00n
MM1 m pm VDD VNW p18 W=0.69u L=180.00n
MM7 pm cn net56 VNW p18 W=0.42u L=180.00n
MM6 net56 m VDD VNW p18 W=0.42u L=180.00n
MM11 net17 m VDD VNW p18 W=2.02u L=180.00n
MM12 net17 c VDD VNW p18 W=2.02u L=180.00n
MM16 Q net17 VDD VNW p18 W=6.06u L=180.00n
MM24 net84 TE VDD VNW p18 W=0.975u L=180.00n
MM0 pm c net80 VNW p18 W=0.975u L=180.00n
MM2 net80 E net84 VNW p18 W=0.975u L=180.00n
MM18 cn CK VDD VNW p18 W=0.88u L=180.00n
MM20 c cn VDD VNW p18 W=800.00n L=180.00n
.ENDS CLKLANQUHDV6
.SUBCKT CLKLANQUHDV8 CK E Q TE VDD VSS VNW VPW
MM4 m pm VSS VPW n18 W=0.47u L=180.00n
MM9 net243 m VSS VPW n18 W=0.43u L=180.00n
MM8 pm c net243 VPW n18 W=0.43u L=180.00n
MM13 net235 c net231 VPW n18 W=1.44u L=180.00n
MM14 net231 m VSS VPW n18 W=1.44u L=180.00n
MM17 Q net235 VSS VPW n18 W=3.25u L=180.00n
MM25 net219 E VSS VPW n18 W=0.47u L=180.00n
MM5 net219 TE VSS VPW n18 W=0.47u L=180.00n
MM3 pm cn net219 VPW n18 W=0.47u L=180.00n
MM19 cn CK VSS VPW n18 W=0.58u L=180.00n
MM21 c cn VSS VPW n18 W=0.58u L=180.00n
MM1 m pm VDD VNW p18 W=0.69u L=180.00n
MM7 pm cn net202 VNW p18 W=0.42u L=180.00n
MM6 net202 m VDD VNW p18 W=0.42u L=180.00n
MM11 net235 m VDD VNW p18 W=2.18u L=180.00n
MM12 net235 c VDD VNW p18 W=2.18u L=180.00n
MM16 Q net235 VDD VNW p18 W=8.6u L=180.00n
MM24 net174 TE VDD VNW p18 W=0.975u L=180.00n
MM0 pm c net178 VNW p18 W=0.975u L=180.00n
MM2 net178 E net174 VNW p18 W=0.975u L=180.00n
MM18 cn CK VDD VNW p18 W=0.88u L=180.00n
MM20 c cn VDD VNW p18 W=0.88u L=180.00n
.ENDS CLKLANQUHDV8
.SUBCKT CLKMUX2UHDV0P7 I0 I1 S Z VDD VSS VNW VPW
MM12 SN S VSS VPW n18 W=430.00n L=180.00n
MM0 net79 SN net75 VPW n18 W=430.00n L=180.00n
MM3 net75 I0 VSS VPW n18 W=430.00n L=180.00n
MM4 net71 I1 VSS VPW n18 W=430.00n L=180.00n
MM5 net79 S net71 VPW n18 W=430.00n L=180.00n
MM8 Z net79 VSS VPW n18 W=430.00n L=180.00n
MM13 SN S VDD VNW p18 W=500.0n L=180.00n
MM1 net79 S net106 VNW p18 W=500.0n L=180.00n
MM2 net106 I0 VDD VNW p18 W=500.0n L=180.00n
MM6 net94 I1 VDD VNW p18 W=500.0n L=180.00n
MM7 net79 SN net94 VNW p18 W=500.0n L=180.00n
MM9 Z net79 VDD VNW p18 W=790.0n L=180.00n
.ENDS CLKMUX2UHDV0P7
.SUBCKT CLKMUX2UHDV1 I0 I1 S Z VDD VSS VNW VPW
MM23 Z net0131 VSS VPW n18 W=430.00n L=180.00n
MM22 net0131 S net0123 VPW n18 W=430.00n L=180.00n
MM21 net0123 I1 VSS VPW n18 W=430.00n L=180.00n
MM20 net0127 I0 VSS VPW n18 W=430.00n L=180.00n
MM19 net0131 SN net0127 VPW n18 W=430.00n L=180.00n
MM18 SN S VSS VPW n18 W=430.00n L=180.00n
MM17 Z net0131 VDD VNW p18 W=1.01u L=180.00n
MM16 net0131 SN net0170 VNW p18 W=0.52u L=180.00n
MM15 net0170 I1 VDD VNW p18 W=0.52u L=180.00n
MM14 net0182 I0 VDD VNW p18 W=0.52u L=180.00n
MM12 net0131 S net0182 VNW p18 W=0.52u L=180.00n
MM13 SN S VDD VNW p18 W=0.52u L=180.00n
.ENDS CLKMUX2UHDV1
.SUBCKT CLKMUX2UHDV2 I0 I1 S Z VDD VSS VNW VPW
MM12 SN S VSS VPW n18 W=430.00n L=180.00n
MM0 net131 SN net127 VPW n18 W=430.00n L=180.00n
MM3 net127 I0 VSS VPW n18 W=430.00n L=180.00n
MM4 net123 I1 VSS VPW n18 W=430.00n L=180.00n
MM5 net131 S net123 VPW n18 W=430.00n L=180.00n
MM8 Z net131 VSS VPW n18 W=0.72u L=180.00n
MM13 SN S VDD VNW p18 W=0.72u L=180.00n
MM1 net131 S net158 VNW p18 W=0.52u L=180.00n
MM2 net158 I0 VDD VNW p18 W=720.0n L=180.00n
MM6 net146 I1 VDD VNW p18 W=1.01u L=180.00n
MM7 net131 SN net146 VNW p18 W=1.01u L=180.00n
MM9 Z net131 VDD VNW p18 W=2.02u L=180.00n
.ENDS CLKMUX2UHDV2
.SUBCKT CLKMUX2UHDV3 I0 I1 S Z VDD VSS VNW VPW
MM12 SN S VSS VPW n18 W=630.00n L=180.00n
MM0 net131 SN net127 VPW n18 W=430.00n L=180.00n
MM4 net123 I1 VSS VPW n18 W=430.00n L=180.00n
MM3 net127 I0 VSS VPW n18 W=430.00n L=180.00n
MM8 Z net131 VSS VPW n18 W=1180.00n L=180.00n
MM5 net131 S net123 VPW n18 W=430.00n L=180.00n
MM13 SN S VDD VNW p18 W=960.0n L=180.00n
MM1 net131 S net158 VNW p18 W=0.52u L=180.00n
MM2 net158 I0 VDD VNW p18 W=800.0n L=180.00n
MM6 net146 I1 VDD VNW p18 W=1.01u L=180.00n
MM7 net131 SN net146 VNW p18 W=1.01u L=180.00n
MM9 Z net131 VDD VNW p18 W=3.03u L=180.00n
.ENDS CLKMUX2UHDV3
.SUBCKT CLKMUX2UHDV4 I0 I1 S Z VDD VSS VNW VPW
MM12 SN S VSS VPW n18 W=630.00n L=180.00n
MM0 net135 SN net131 VPW n18 W=430.00n L=180.00n
MM3 net131 I0 VSS VPW n18 W=430.00n L=180.00n
MM4 net127 I1 VSS VPW n18 W=430.00n L=180.00n
MM5 net135 S net127 VPW n18 W=430.00n L=180.00n
MM8 Z net135 VSS VPW n18 W=1.58u L=180.00n
MM1 net135 S net162 VNW p18 W=1.305u L=180.00n
MM2 net162 I0 VDD VNW p18 W=1.005u L=180.00n
MM6 net150 I1 VDD VNW p18 W=1.305u L=180.00n
MM7 net135 SN net150 VNW p18 W=1.305u L=180.00n
MM9 Z net135 VDD VNW p18 W=4.04u L=180.00n
MM13 SN S VDD VNW p18 W=960.0n L=180.00n
.ENDS CLKMUX2UHDV4
.SUBCKT CLKMUX2UHDV6 I0 I1 S Z VDD VSS VNW VPW
MM0 net83 SN net79 VPW n18 W=640.00n L=180.00n
MM3 net79 I0 VSS VPW n18 W=640.00n L=180.00n
MM4 net75 I1 VSS VPW n18 W=640.00n L=180.00n
MM5 net83 S net75 VPW n18 W=640.00n L=180.00n
MM8 Z net83 VSS VPW n18 W=2.52u L=180.00n
MM12 SN S VSS VPW n18 W=960.00n L=180.00n
MM1 net83 S net110 VNW p18 W=2.02u L=180.00n
MM2 net110 I0 VDD VNW p18 W=2.02u L=180.00n
MM6 net98 I1 VDD VNW p18 W=2.12u L=180.00n
MM7 net83 SN net98 VNW p18 W=2.12u L=180.00n
MM9 Z net83 VDD VNW p18 W=6.115u L=180.00n
MM13 SN S VDD VNW p18 W=1.45u L=180.00n
.ENDS CLKMUX2UHDV6
.SUBCKT CLKMUX2UHDV8 I0 I1 S Z VDD VSS VNW VPW
MM12 SN S VSS VPW n18 W=1.35u L=180.00n
MM0 net135 SN net131 VPW n18 W=1030.00n L=180.00n
MM3 net131 I0 VSS VPW n18 W=1030.00n L=180.00n
MM4 net127 I1 VSS VPW n18 W=1030.00n L=180.00n
MM5 net135 S net127 VPW n18 W=1030.00n L=180.00n
MM8 Z net135 VSS VPW n18 W=3.16u L=180.00n
MM1 net135 S net162 VNW p18 W=2.85u L=180.00n
MM2 net162 I0 VDD VNW p18 W=3.03u L=180.00n
MM6 net150 I1 VDD VNW p18 W=3.27u L=180.00n
MM7 net135 SN net150 VNW p18 W=2.85u L=180.00n
MM9 Z net135 VDD VNW p18 W=8.57u L=180.00n
MM13 SN S VDD VNW p18 W=2.19u L=180.00n
.ENDS CLKMUX2UHDV8
.SUBCKT CLKNAND2UHDV0P7 A1 A2 ZN VDD VSS VNW VPW
MM3 ZN A1 net16 VPW n18 W=370.00n L=180.00n
MM5 net16 A2 VSS VPW n18 W=370.00n L=180.00n
MM2 ZN A1 VDD VNW p18 W=710.0n L=180.00n
MM0 ZN A2 VDD VNW p18 W=710.0n L=180.00n
.ENDS CLKNAND2UHDV0P7
.SUBCKT CLKNAND2UHDV1 A1 A2 ZN VDD VSS VNW VPW
MM5 net4 A2 VSS VPW n18 W=530.00n L=180.00n
MM3 ZN A1 net4 VPW n18 W=530.00n L=180.00n
MM0 ZN A2 VDD VNW p18 W=1.01u L=180.00n
MM2 ZN A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKNAND2UHDV1
.SUBCKT CLKNAND2UHDV2 A1 A2 ZN VDD VSS VNW VPW
MM3 ZN A1 net16 VPW n18 W=1.06u L=180.00n
MM5 net16 A2 VSS VPW n18 W=1.06u L=180.00n
MM2 ZN A1 VDD VNW p18 W=1.9u L=180.00n
MM0 ZN A2 VDD VNW p18 W=2.02u L=180.00n
.ENDS CLKNAND2UHDV2
.SUBCKT CLKNAND2UHDV3 A1 A2 ZN VDD VSS VNW VPW
MM5 net4 A2 VSS VPW n18 W=1.59u L=180.00n
MM3 ZN A1 net4 VPW n18 W=1.59u L=180.00n
MM0 ZN A2 VDD VNW p18 W=2.97u L=180.00n
MM2 ZN A1 VDD VNW p18 W=2.85u L=180.00n
.ENDS CLKNAND2UHDV3
.SUBCKT CLKNAND2UHDV4 A1 A2 ZN VDD VSS VNW VPW
MM5 net4 A2 VSS VPW n18 W=2.12u L=180.00n
MM3 ZN A1 net4 VPW n18 W=2.12u L=180.00n
MM0 ZN A2 VDD VNW p18 W=3.98u L=180.00n
MM2 ZN A1 VDD VNW p18 W=3.86u L=180.00n
.ENDS CLKNAND2UHDV4
.SUBCKT CLKNAND2UHDV6 A1 A2 ZN VDD VSS VNW VPW
MM3 ZN A1 net16 VPW n18 W=3.18u L=180.00n
MM5 net16 A2 VSS VPW n18 W=3.18u L=180.00n
MM2 ZN A1 VDD VNW p18 W=4.75u L=180.00n
MM0 ZN A2 VDD VNW p18 W=4.99u L=180.00n
.ENDS CLKNAND2UHDV6
.SUBCKT CLKNAND2UHDV8 A1 A2 ZN VDD VSS VNW VPW
MM3 ZN A1 net16 VPW n18 W=4.24u L=180.00n
MM5 net16 A2 VSS VPW n18 W=4.24u L=180.00n
MM2 ZN A1 VDD VNW p18 W=7.66u L=180.00n
MM0 ZN A2 VDD VNW p18 W=8.08u L=180.00n
.ENDS CLKNAND2UHDV8
.SUBCKT CLKNOR2UHDV0P7 A1 A2 ZN VDD VSS VNW VPW
MM5 ZN A2 VSS VPW n18 W=250.00n L=180.00n
MM9 ZN A1 VSS VPW n18 W=250.00n L=180.00n
MM4 net19 A2 VDD VNW p18 W=710.0n L=180.00n
MM8 ZN A1 net19 VNW p18 W=710.0n L=180.00n
.ENDS CLKNOR2UHDV0P7
.SUBCKT CLKNOR2UHDV1 A1 A2 ZN VDD VSS VNW VPW
MM9 ZN A1 VSS VPW n18 W=250.00n L=180.00n
MM5 ZN A2 VSS VPW n18 W=250.00n L=180.00n
MM8 ZN A1 net7 VNW p18 W=1.01u L=180.00n
MM4 net7 A2 VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKNOR2UHDV1
.SUBCKT CLKNOR2UHDV2 A1 A2 ZN VDD VSS VNW VPW
MM9 ZN A1 VSS VPW n18 W=500.00n L=180.00n
MM5 ZN A2 VSS VPW n18 W=500.00n L=180.00n
MM8 ZN A1 net7 VNW p18 W=2.02u L=180.00n
MM4 net7 A2 VDD VNW p18 W=2.02u L=180.00n
.ENDS CLKNOR2UHDV2
.SUBCKT CLKNOR2UHDV3 A1 A2 ZN VDD VSS VNW VPW
MM9 ZN A1 VSS VPW n18 W=750.00n L=180.00n
MM5 ZN A2 VSS VPW n18 W=750.00n L=180.00n
MM8 ZN A1 net7 VNW p18 W=3.03u L=180.00n
MM4 net7 A2 VDD VNW p18 W=3.03u L=180.00n
.ENDS CLKNOR2UHDV3
.SUBCKT CLKNOR2UHDV4 A1 A2 ZN VDD VSS VNW VPW
MM9 ZN A1 VSS VPW n18 W=1u L=180.00n
MM5 ZN A2 VSS VPW n18 W=1u L=180.00n
MM8 ZN A1 net7 VNW p18 W=4.04u L=180.00n
MM4 net7 A2 VDD VNW p18 W=4.04u L=180.00n
.ENDS CLKNOR2UHDV4
.SUBCKT CLKNOR2UHDV6 A1 A2 ZN VDD VSS VNW VPW
MM9 ZN A1 VSS VPW n18 W=1.5u L=180.00n
MM5 ZN A2 VSS VPW n18 W=1.5u L=180.00n
MM8 ZN A1 net7 VNW p18 W=6.06u L=180.00n
MM4 net7 A2 VDD VNW p18 W=6.06u L=180.00n
.ENDS CLKNOR2UHDV6
.SUBCKT CLKNOR2UHDV8 A1 A2 ZN VDD VSS VNW VPW
MM9 ZN A1 VSS VPW n18 W=2u L=180.00n
MM5 ZN A2 VSS VPW n18 W=2u L=180.00n
MM8 ZN A1 net7 VNW p18 W=8.48u L=180.00n
MM4 net7 A2 VDD VNW p18 W=8.48u L=180.00n
.ENDS CLKNOR2UHDV8
.SUBCKT CLKOR2UHDV0P7 A1 A2 Z VDD VSS VNW VPW
MM6 Z net20 VDD VNW p18 W=790.00n L=180.00n
MM7 net15 A2 VDD VNW p18 W=500.00n L=180.00n
MM0 net20 A1 net15 VNW p18 W=500.00n L=180.00n
MM8 Z net20 VSS VPW n18 W=430.00n L=180.00n
MM15 net20 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 net20 A1 VSS VPW n18 W=430.00n L=180.00n
.ENDS CLKOR2UHDV0P7
.SUBCKT CLKOR2UHDV1 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=430.00n L=180.00n
MM15 net8 A2 VSS VPW n18 W=430.00n L=180.00n
MM8 Z net8 VSS VPW n18 W=430.00n L=180.00n
MM0 net8 A1 net19 VNW p18 W=810.00n L=180.00n
MM7 net19 A2 VDD VNW p18 W=810.00n L=180.00n
MM6 Z net8 VDD VNW p18 W=1.01u L=180.00n
.ENDS CLKOR2UHDV1
.SUBCKT CLKOR2UHDV2 A1 A2 Z VDD VSS VNW VPW
MM6 Z net20 VDD VNW p18 W=2.02u L=180.00n
MM7 net15 A2 VDD VNW p18 W=1.01u L=180.00n
MM0 net20 A1 net15 VNW p18 W=1.01u L=180.00n
MM8 Z net20 VSS VPW n18 W=1.18u L=180.00n
MM15 net20 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 net20 A1 VSS VPW n18 W=430.00n L=180.00n
.ENDS CLKOR2UHDV2
.SUBCKT CLKOR2UHDV3 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=430.00n L=180.00n
MM15 net8 A2 VSS VPW n18 W=430.00n L=180.00n
MM8 Z net8 VSS VPW n18 W=1180.00n L=180.00n
MM0 net8 A1 net19 VNW p18 W=1.01u L=180.00n
MM7 net19 A2 VDD VNW p18 W=1.01u L=180.00n
MM6 Z net8 VDD VNW p18 W=3.03u L=180.00n
.ENDS CLKOR2UHDV3
.SUBCKT CLKOR2UHDV4 A1 A2 Z VDD VSS VNW VPW
MM6 Z net20 VDD VNW p18 W=4.04u L=180.00n
MM7 net15 A2 VDD VNW p18 W=1.355u L=180.00n
MM0 net20 A1 net15 VNW p18 W=1.41u L=180.00n
MM8 Z net20 VSS VPW n18 W=1.57u L=180.00n
MM15 net20 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 net20 A1 VSS VPW n18 W=430.00n L=180.00n
.ENDS CLKOR2UHDV4
.SUBCKT CLKOR2UHDV6 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=640.00n L=180.00n
MM15 net8 A2 VSS VPW n18 W=640.00n L=180.00n
MM8 Z net8 VSS VPW n18 W=2.38u L=180.00n
MM0 net8 A1 net19 VNW p18 W=1.96u L=180.00n
MM7 net19 A2 VDD VNW p18 W=1.96u L=180.00n
MM6 Z net8 VDD VNW p18 W=5.88u L=180.00n
.ENDS CLKOR2UHDV6
.SUBCKT CLKOR2UHDV8 A1 A2 Z VDD VSS VNW VPW
MM6 Z net20 VDD VNW p18 W=8.39u L=180.00n
MM7 net15 A2 VDD VNW p18 W=3.36u L=180.00n
MM0 net20 A1 net15 VNW p18 W=3.26u L=180.00n
MM8 Z net20 VSS VPW n18 W=3.12u L=180.00n
MM15 net20 A2 VSS VPW n18 W=1.04u L=180.00n
MM3 net20 A1 VSS VPW n18 W=1030.00n L=180.00n
.ENDS CLKOR2UHDV8
.SUBCKT CLKXOR2UHDV0P7 A1 A2 Z VDD VSS VNW VPW
MM6 Z A1 net7 VNW p18 W=790.0n L=180.00n
MM5 net7 a2n VDD VNW p18 W=790.0n L=180.00n
MM11 a2n a1n Z VNW p18 W=790.0n L=180.00n
MM2 a1n A1 VDD VNW p18 W=790.0n L=180.00n
MM1 a2n A2 VDD VNW p18 W=790.0n L=180.00n
MM7 Z a1n net28 VPW n18 W=430.00n L=180.00n
MM4 net28 a2n VSS VPW n18 W=430.00n L=180.00n
MM13 a2n A1 Z VPW n18 W=430.00n L=180.00n
MM3 a1n A1 VSS VPW n18 W=430.00n L=180.00n
MM0 a2n A2 VSS VPW n18 W=430.00n L=180.00n
.ENDS CLKXOR2UHDV0P7
.SUBCKT CLKXOR2UHDV1 A1 A2 Z VDD VSS VNW VPW
MM6 Z A1 net7 VNW p18 W=1.01u L=180.00n
MM5 net7 a2n VDD VNW p18 W=1.01u L=180.00n
MM11 a2n a1n Z VNW p18 W=1.01u L=180.00n
MM2 a1n A1 VDD VNW p18 W=1.01u L=180.00n
MM1 a2n A2 VDD VNW p18 W=1.01u L=180.00n
MM0 a2n A2 VSS VPW n18 W=430.00n L=180.00n
MM7 Z a1n net32 VPW n18 W=430.00n L=180.00n
MM4 net32 a2n VSS VPW n18 W=430.00n L=180.00n
MM13 a2n A1 Z VPW n18 W=430.00n L=180.00n
MM3 a1n A1 VSS VPW n18 W=430.00n L=180.00n
.ENDS CLKXOR2UHDV1
.SUBCKT CLKXOR2UHDV2 A1 A2 Z VDD VSS VNW VPW
MM0 a2n A2 VSS VPW n18 W=0.86u L=180.00n
MM3 a1n A1 VSS VPW n18 W=0.84u L=180.00n
MM13 a2n A1 Z VPW n18 W=720.00n L=180.00n
MM8 net20 a1n Z VPW n18 W=0.825u L=180.00n
MM9 net20 a2n VSS VPW n18 W=430.00n L=180.00n
MM1 a2n A2 VDD VNW p18 W=2.02u L=180.00n
MM2 a1n A1 VDD VNW p18 W=2.02u L=180.00n
MM11 a2n a1n Z VNW p18 W=0.925u L=180.00n
MM7 net20 A1 Z VNW p18 W=0.925u L=180.00n
MM10 net20 a2n VDD VNW p18 W=0.925u L=180.00n
.ENDS CLKXOR2UHDV2
.SUBCKT CLKXOR2UHDV4 A1 A2 Z VDD VSS VNW VPW
MM9 net4 a2n VSS VPW n18 W=430.00n L=180.00n
MM8 net4 a1n Z VPW n18 W=2.23u L=180.00n
MM13 a2n A1 Z VPW n18 W=2.33u L=180.00n
MM3 a1n A1 VSS VPW n18 W=1.58u L=180.00n
MM0 a2n A2 VSS VPW n18 W=1.58u L=180.00n
MM10 net4 a2n VDD VNW p18 W=1.01u L=180.00n
MM7 net4 A1 Z VNW p18 W=2.775u L=180.00n
MM11 a2n a1n Z VNW p18 W=3.35u L=180.00n
MM2 a1n A1 VDD VNW p18 W=4.04u L=180.00n
MM1 a2n A2 VDD VNW p18 W=4.04u L=180.00n
.ENDS CLKXOR2UHDV4
****Sub-Circuit for DEL1UHDV1, Fri Nov  6 11:29:59 CST 2015****
.SUBCKT DEL1UHDV1 I Z VDD VSS VNW VPW
MM6 net044 I VDD VNW p18 W=350.0n L=180.00n
MM3 net19 net042 VDD VNW p18 W=750.00n L=180.00n
MM1 Z net19 VDD VNW p18 W=1.01u L=180.00n
MM4 net042 net044 VDD VNW p18 W=750.00n L=180.00n
MM7 net044 I VSS VPW n18 W=250.00n L=180.00n
MM2 net19 net042 VSS VPW n18 W=250.00n L=180.00n
MM0 Z net19 VSS VPW n18 W=320.00n L=180.00n
MM5 net042 net044 VSS VPW n18 W=250.00n L=180.00n
.ENDS DEL1UHDV1
****Sub-Circuit for DEL1UHDV2, Fri Nov  6 11:29:59 CST 2015****
.SUBCKT DEL1UHDV2 I Z VDD VSS VNW VPW
MM6 net044 I VDD VNW p18 W=370.0n L=180.00n
MM3 net19 net042 VDD VNW p18 W=850.00n L=180.00n
MM1 Z net19 VDD VNW p18 W=2.02u L=180.00n
MM4 net042 net044 VDD VNW p18 W=850.00n L=180.00n
MM7 net044 I VSS VPW n18 W=250.00n L=180.00n
MM2 net19 net042 VSS VPW n18 W=250.00n L=180.00n
MM0 Z net19 VSS VPW n18 W=730.00n L=180.00n
MM5 net042 net044 VSS VPW n18 W=250.00n L=180.00n
.ENDS DEL1UHDV2
****Sub-Circuit for DEL2UHDV1, Fri Nov  6 11:29:59 CST 2015****
.SUBCKT DEL2UHDV1 I Z VDD VSS VNW VPW
MM4 net029 net046 VDD VNW p18 W=840.00n L=180.00n
MM5 net050 net046 net029 VNW p18 W=840.00n L=180.00n
MM9 net046 I VDD VNW p18 W=700n L=180.00n
MM3 net10 net050 VDD VNW p18 W=840.00n L=180.00n
MM7 net19 net050 net10 VNW p18 W=840.00n L=180.00n
MM1 Z net19 VDD VNW p18 W=1.01u L=180.00n
MM6 net054 net046 VSS VPW n18 W=250.00n L=180.00n
MM8 net050 net046 net054 VPW n18 W=250.00n L=180.00n
MM10 net046 I VSS VPW n18 W=250.00n L=180.00n
MM2 net15 net050 VSS VPW n18 W=250.00n L=180.00n
MM15 net19 net050 net15 VPW n18 W=250.00n L=180.00n
MM0 Z net19 VSS VPW n18 W=360.00n L=180.00n
.ENDS DEL2UHDV1
****Sub-Circuit for DEL2UHDV2, Fri Nov  6 11:29:59 CST 2015****
.SUBCKT DEL2UHDV2 I Z VDD VSS VNW VPW
MM7 net19 net058 net029 VNW p18 W=900.00n L=180.00n
MM11 net029 net058 VDD VNW p18 W=900.00n L=180.00n
MM9 net054 I VDD VNW p18 W=720n L=180.00n
MM4 net037 net054 VDD VNW p18 W=900.00n L=180.00n
MM1 Z net19 VDD VNW p18 W=2.02u L=180.00n
MM5 net058 net054 net037 VNW p18 W=900.00n L=180.00n
MM3 net19 net058 net046 VPW n18 W=250.00n L=180.00n
MM12 net046 net058 VSS VPW n18 W=250.00n L=180.00n
MM6 net062 net054 VSS VPW n18 W=250.00n L=180.00n
MM8 net058 net054 net062 VPW n18 W=250.00n L=180.00n
MM0 Z net19 VSS VPW n18 W=720.00n L=180.00n
MM10 net054 I VSS VPW n18 W=250.00n L=180.00n
.ENDS DEL2UHDV2
****Sub-Circuit for DEL4UHDV1, Fri Nov  6 11:29:59 CST 2015****
.SUBCKT DEL4UHDV1 I Z VDD VSS VNW VPW
MM13 net057 I VDD VNW p18 W=490.00n L=180.00n
MM4 net036 net057 net051 VNW p18 W=840.00n L=180.00n
MM5 net061 net057 net036 VNW p18 W=840.00n L=180.00n
MM14 net063 net057 VDD VNW p18 W=840.00n L=180.00n
MM16 net051 net057 net063 VNW p18 W=840.00n L=180.00n
MM17 net071 net061 VDD VNW p18 W=840.00n L=180.00n
MM18 net075 net061 net071 VNW p18 W=840.00n L=180.00n
MM3 net10 net061 net075 VNW p18 W=840.00n L=180.00n
MM7 net19 net061 net10 VNW p18 W=840.00n L=180.00n
MM1 Z net19 VDD VNW p18 W=1.01u L=180.00n
MM20 net088 net061 VSS VPW n18 W=250.00n L=180.00n
MM21 net084 net061 net088 VPW n18 W=250.00n L=180.00n
MM11 net057 I VSS VPW n18 W=250.00n L=180.00n
MM6 net065 net057 net092 VPW n18 W=250.00n L=180.00n
MM8 net061 net057 net065 VPW n18 W=250.00n L=180.00n
MM12 net096 net057 VSS VPW n18 W=250.00n L=180.00n
MM19 net092 net057 net096 VPW n18 W=250.00n L=180.00n
MM2 net15 net061 net084 VPW n18 W=250.00n L=180.00n
MM15 net19 net061 net15 VPW n18 W=250.00n L=180.00n
MM0 Z net19 VSS VPW n18 W=340.00n L=180.00n
.ENDS DEL4UHDV1
****Sub-Circuit for DEL4UHDV2, Fri Nov  6 11:29:59 CST 2015****
.SUBCKT DEL4UHDV2 I Z VDD VSS VNW VPW
MM37 net064 net052 VSS VPW n18 W=250.00n L=180.00n
MM38 net060 net052 net056 VPW n18 W=250.00n L=180.00n
MM39 net056 net052 net068 VPW n18 W=250.00n L=180.00n
MM51 net052 I VSS VPW n18 W=250.00n L=180.00n
MM41 net048 net060 net044 VPW n18 W=250.00n L=180.00n
MM42 net044 net060 VSS VPW n18 W=250.00n L=180.00n
MM34 net111 net060 net072 VPW n18 W=250.00n L=180.00n
MM35 net072 net060 net048 VPW n18 W=250.00n L=180.00n
MM36 net068 net052 net064 VPW n18 W=250.00n L=180.00n
MM0 Z net111 VSS VPW n18 W=840.00n L=180.00n
MM52 net052 I VDD VNW p18 W=490.00n L=180.00n
MM43 net111 net060 net0119 VNW p18 W=910.00n L=180.00n
MM44 net0119 net060 net0115 VNW p18 W=910.00n L=180.00n
MM45 net0115 net060 net0111 VNW p18 W=910.00n L=180.00n
MM46 net0111 net060 VDD VNW p18 W=910.00n L=180.00n
MM47 net091 net052 net0103 VNW p18 W=910.00n L=180.00n
MM48 net0103 net052 VDD VNW p18 W=910.00n L=180.00n
MM49 net060 net052 net095 VNW p18 W=910.00n L=180.00n
MM50 net095 net052 net091 VNW p18 W=910.00n L=180.00n
MM1 Z net111 VDD VNW p18 W=2.02u L=180.00n
.ENDS DEL4UHDV2
****Sub-Circuit for DGRNQNUHDV0P7, Thu Jun  8 09:36:16 CST 2017****
.SUBCKT DGRNQNUHDV0P7 CK D QN RN VDD VSS VNW VPW
MM31 net0136 cn net83 VPW n18 W=0.5u L=180.00n
MM20 net0132 net83 VSS VPW n18 W=0.5u L=180.00n
MM18 net0136 net0132 VSS VPW n18 W=0.5u L=180.00n
MM16 net0112 c net83 VPW n18 W=0.43u L=180.00n
MM15 net0120 net0112 VSS VPW n18 W=0.36u L=180.00n
MM13 net0111 c net0120 VPW n18 W=0.73u L=180.00n
MM10 net0112 net0111 VSS VPW n18 W=0.36u L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM7 net0102 D net094 VPW n18 W=360.00n L=180.00n
MM9 net0111 cn net0102 VPW n18 W=360.00n L=180.00n
MM38 net094 RN VSS VPW n18 W=360.00n L=180.00n
MM24 QN net83 VSS VPW n18 W=560.00n L=180.00n
MM8 net0146 D VDD VNW p18 W=580.00n L=180.00n
MM4 net0111 c net0146 VNW p18 W=580.00n L=180.00n
MM37 net0146 RN VDD VNW p18 W=580.00n L=180.00n
MM23 net0132 net83 VDD VNW p18 W=1.01u L=180.00n
MM22 net0176 net0132 VDD VNW p18 W=0.73u L=180.00n
MM26 net0176 c net83 VNW p18 W=0.49u L=180.00n
MM17 net0112 cn net83 VNW p18 W=820.00n L=180.00n
MM14 net0111 cn net0171 VNW p18 W=580.00n L=180.00n
MM12 net0171 net0112 VDD VNW p18 W=0.58u L=180.00n
MM11 net0112 net0111 VDD VNW p18 W=450.00n L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM25 QN net83 VDD VNW p18 W=810.0n L=180.00n
.ENDS DGRNQNUHDV0P7
****Sub-Circuit for DGRNQNUHDV1, Thu Jun  8 09:36:16 CST 2017****
.SUBCKT DGRNQNUHDV1 CK D QN RN VDD VSS VNW VPW
MM10 net0132 net0139 VSS VPW n18 W=0.36u L=180.00n
MM13 net0139 c net0124 VPW n18 W=0.73u L=180.00n
MM15 net0124 net0132 VSS VPW n18 W=0.36u L=180.00n
MM31 net0120 cn net23 VPW n18 W=0.5u L=180.00n
MM16 net0132 c net23 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM20 net0100 net23 VSS VPW n18 W=0.5u L=180.00n
MM18 net0120 net0100 VSS VPW n18 W=0.5u L=180.00n
MM7 net0102 D net094 VPW n18 W=360.00n L=180.00n
MM9 net0139 cn net0102 VPW n18 W=360.00n L=180.00n
MM38 net094 RN VSS VPW n18 W=360.00n L=180.00n
MM24 QN net23 VSS VPW n18 W=720.00n L=180.00n
MM11 net0132 net0139 VDD VNW p18 W=450.00n L=180.00n
MM12 net0175 net0132 VDD VNW p18 W=0.58u L=180.00n
MM14 net0139 cn net0175 VNW p18 W=580.00n L=180.00n
MM26 net0168 c net23 VNW p18 W=0.49u L=180.00n
MM17 net0132 cn net23 VNW p18 W=820.00n L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM23 net0100 net23 VDD VNW p18 W=1.01u L=180.00n
MM22 net0168 net0100 VDD VNW p18 W=0.73u L=180.00n
MM8 net0146 D VDD VNW p18 W=580.00n L=180.00n
MM4 net0139 c net0146 VNW p18 W=580.00n L=180.00n
MM37 net0146 RN VDD VNW p18 W=580.00n L=180.00n
MM25 QN net23 VDD VNW p18 W=1.01u L=180.00n
.ENDS DGRNQNUHDV1
****Sub-Circuit for DGRNQNUHDV2, Thu Jun  8 09:36:16 CST 2017****
.SUBCKT DGRNQNUHDV2 CK D QN RN VDD VSS VNW VPW
MM9 net187 cn net0109 VPW n18 W=360.00n L=180.00n
MM38 net0101 RN VSS VPW n18 W=360.00n L=180.00n
MM10 net180 net187 VSS VPW n18 W=0.34u L=180.00n
MM13 net187 c net172 VPW n18 W=0.73u L=180.00n
MM15 net172 net180 VSS VPW n18 W=0.34u L=180.00n
MM31 net168 cn net167 VPW n18 W=0.53u L=180.00n
MM20 net148 net167 VSS VPW n18 W=0.53u L=180.00n
MM18 net168 net148 VSS VPW n18 W=0.53u L=180.00n
MM16 net180 c net167 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM24 QN net167 VSS VPW n18 W=1.44u L=180.00n
MM7 net0109 D net0101 VPW n18 W=360.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM12 net127 net180 VDD VNW p18 W=580.00n L=180.00n
MM14 net187 cn net127 VNW p18 W=580.00n L=180.00n
MM26 net120 c net167 VNW p18 W=0.49u L=180.00n
MM17 net180 cn net167 VNW p18 W=820.00n L=180.00n
MM11 net180 net187 VDD VNW p18 W=450.00n L=180.00n
MM23 net148 net167 VDD VNW p18 W=1.01u L=180.00n
MM8 net0153 D VDD VNW p18 W=580.00n L=180.00n
MM4 net187 c net0153 VNW p18 W=580.00n L=180.00n
MM37 net0153 RN VDD VNW p18 W=580.00n L=180.00n
MM22 net120 net148 VDD VNW p18 W=0.73u L=180.00n
MM25 QN net167 VDD VNW p18 W=2.02u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
.ENDS DGRNQNUHDV2
****Sub-Circuit for DGRSNQNUHDV0P7, Mon Jun 26 14:26:51 CST 2017****
.SUBCKT DGRSNQNUHDV0P7 CK D QN RN SN VDD VSS VNW VPW
MM5 snn SN VSS VPW n18 W=280.00n L=180.00n
MM42 net0122 snn net0114 VPW n18 W=420.00n L=180.00n
MM31 net0136 cn net83 VPW n18 W=0.5u L=180.00n
MM20 net0132 net83 VSS VPW n18 W=420.00n L=180.00n
MM38 net0114 RN VSS VPW n18 W=420.00n L=180.00n
MM9 net0111 cn net0122 VPW n18 W=430.00n L=180.00n
MM7 net0122 D net0114 VPW n18 W=420.00n L=180.00n
MM18 net0136 net0132 VSS VPW n18 W=0.5u L=180.00n
MM16 net0112 c net83 VPW n18 W=0.43u L=180.00n
MM15 net0120 net0112 VSS VPW n18 W=430.00n L=180.00n
MM13 net0111 c net0120 VPW n18 W=430.00n L=180.00n
MM10 net0112 net0111 VSS VPW n18 W=0.36u L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM24 QN net83 VSS VPW n18 W=560.00n L=180.00n
MM6 snn SN VDD VNW p18 W=420.00n L=180.00n
MM41 net0109 snn VDD VNW p18 W=580.00n L=180.00n
MM37 net098 RN VDD VNW p18 W=580.00n L=180.00n
MM4 net0111 c net098 VNW p18 W=580.00n L=180.00n
MM8 net098 D net0109 VNW p18 W=580.00n L=180.00n
MM23 net0132 net83 VDD VNW p18 W=420.00n L=180.00n
MM22 net0176 net0132 VDD VNW p18 W=490.00n L=180.00n
MM26 net0176 c net83 VNW p18 W=0.49u L=180.00n
MM17 net0112 cn net83 VNW p18 W=565.00n L=180.00n
MM14 net0111 cn net0171 VNW p18 W=580.00n L=180.00n
MM12 net0171 net0112 VDD VNW p18 W=0.58u L=180.00n
MM11 net0112 net0111 VDD VNW p18 W=0.58u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM25 QN net83 VDD VNW p18 W=810.0n L=180.00n
.ENDS DGRSNQNUHDV0P7
****Sub-Circuit for DGRSNQNUHDV1, Mon Jun 26 14:26:51 CST 2017****
.SUBCKT DGRSNQNUHDV1 CK D QN RN SN VDD VSS VNW VPW
MM5 snn SN VSS VPW n18 W=280.00n L=180.00n
MM10 net0132 net0139 VSS VPW n18 W=0.36u L=180.00n
MM13 net0139 c net0124 VPW n18 W=430.00n L=180.00n
MM15 net0124 net0132 VSS VPW n18 W=430.00n L=180.00n
MM31 net0120 cn net23 VPW n18 W=0.5u L=180.00n
MM16 net0132 c net23 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM20 net0100 net23 VSS VPW n18 W=420.00n L=180.00n
MM18 net0120 net0100 VSS VPW n18 W=0.5u L=180.00n
MM38 net0101 RN VSS VPW n18 W=420.00n L=180.00n
MM42 net098 snn net0101 VPW n18 W=420.00n L=180.00n
MM7 net098 D net0101 VPW n18 W=420.00n L=180.00n
MM9 net0139 cn net098 VPW n18 W=430.00n L=180.00n
MM24 QN net23 VSS VPW n18 W=720.00n L=180.00n
MM6 snn SN VDD VNW p18 W=420.00n L=180.00n
MM11 net0132 net0139 VDD VNW p18 W=0.58u L=180.00n
MM12 net0175 net0132 VDD VNW p18 W=0.58u L=180.00n
MM14 net0139 cn net0175 VNW p18 W=580.00n L=180.00n
MM26 net0168 c net23 VNW p18 W=0.49u L=180.00n
MM17 net0132 cn net23 VNW p18 W=565.00n L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM23 net0100 net23 VDD VNW p18 W=420.00n L=180.00n
MM22 net0168 net0100 VDD VNW p18 W=490.00n L=180.00n
MM4 net0139 c net0150 VNW p18 W=580.00n L=180.00n
MM8 net0150 D net0161 VNW p18 W=580.00n L=180.00n
MM41 net0161 snn VDD VNW p18 W=580.00n L=180.00n
MM37 net0150 RN VDD VNW p18 W=580.00n L=180.00n
MM25 QN net23 VDD VNW p18 W=1.01u L=180.00n
.ENDS DGRSNQNUHDV1
****Sub-Circuit for DGRSNQNUHDV2, Mon Jun 26 14:26:51 CST 2017****
.SUBCKT DGRSNQNUHDV2 CK D QN RN SN VDD VSS VNW VPW
MM5 snn SN VSS VPW n18 W=280.00n L=180.00n
MM9 net187 cn net0101 VPW n18 W=430.00n L=180.00n
MM7 net0101 D net0104 VPW n18 W=420.00n L=180.00n
MM10 net180 net187 VSS VPW n18 W=360.00n L=180.00n
MM13 net187 c net172 VPW n18 W=430.00n L=180.00n
MM15 net172 net180 VSS VPW n18 W=430.00n L=180.00n
MM31 net168 cn net167 VPW n18 W=500.00n L=180.00n
MM20 net148 net167 VSS VPW n18 W=420.00n L=180.00n
MM18 net168 net148 VSS VPW n18 W=500.00n L=180.00n
MM16 net180 c net167 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM42 net0101 snn net0104 VPW n18 W=420.00n L=180.00n
MM38 net0104 RN VSS VPW n18 W=420.00n L=180.00n
MM24 QN net167 VSS VPW n18 W=1.44u L=180.00n
MM6 snn SN VDD VNW p18 W=420.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM12 net127 net180 VDD VNW p18 W=580.00n L=180.00n
MM14 net187 cn net127 VNW p18 W=580.00n L=180.00n
MM26 net120 c net167 VNW p18 W=0.49u L=180.00n
MM17 net180 cn net167 VNW p18 W=565.00n L=180.00n
MM11 net180 net187 VDD VNW p18 W=580.00n L=180.00n
MM23 net148 net167 VDD VNW p18 W=420.00n L=180.00n
MM37 net0161 RN VDD VNW p18 W=580.00n L=180.00n
MM41 net0156 snn VDD VNW p18 W=580.00n L=180.00n
MM8 net0161 D net0156 VNW p18 W=580.00n L=180.00n
MM4 net187 c net0161 VNW p18 W=580.00n L=180.00n
MM22 net120 net148 VDD VNW p18 W=490.00n L=180.00n
MM25 QN net167 VDD VNW p18 W=2.02u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
.ENDS DGRSNQNUHDV2
.SUBCKT DQNUHDV0P7 CK D QN VDD VSS VNW VPW
MM31 net0136 cn net83 VPW n18 W=0.5u L=180.00n
MM20 net0132 net83 VSS VPW n18 W=0.5u L=180.00n
MM18 net0136 net0132 VSS VPW n18 W=0.5u L=180.00n
MM16 net0112 c net83 VPW n18 W=0.43u L=180.00n
MM15 net0120 net0112 VSS VPW n18 W=0.36u L=180.00n
MM13 net0111 c net0120 VPW n18 W=0.73u L=180.00n
MM10 net0112 net0111 VSS VPW n18 W=0.36u L=180.00n
MM9 net096 cn net0111 VPW n18 W=0.5u L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM4 net096 D VSS VPW n18 W=0.36u L=180.00n
MM24 QN net83 VSS VPW n18 W=560.00n L=180.00n
MM23 net0132 net83 VDD VNW p18 W=1.09u L=180.00n
MM22 net0176 net0132 VDD VNW p18 W=0.73u L=180.00n
MM26 net0176 c net83 VNW p18 W=0.49u L=180.00n
MM17 net0112 cn net83 VNW p18 W=0.96u L=180.00n
MM14 net0111 cn net0171 VNW p18 W=580.00n L=180.00n
MM12 net0171 net0112 VDD VNW p18 W=0.58u L=180.00n
MM11 net0112 net0111 VDD VNW p18 W=0.58u L=180.00n
MM6 net0148 c net0111 VNW p18 W=0.58u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM5 net0148 D VDD VNW p18 W=0.58u L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM25 QN net83 VDD VNW p18 W=810.0n L=180.00n
.ENDS DQNUHDV0P7
.SUBCKT DQNUHDV1 CK D QN VDD VSS VNW VPW
MM9 net0104 cn net0139 VPW n18 W=0.5u L=180.00n
MM10 net0132 net0139 VSS VPW n18 W=0.36u L=180.00n
MM13 net0139 c net0124 VPW n18 W=0.73u L=180.00n
MM15 net0124 net0132 VSS VPW n18 W=0.36u L=180.00n
MM31 net0120 cn net23 VPW n18 W=0.5u L=180.00n
MM16 net0132 c net23 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM4 net0104 D VSS VPW n18 W=0.36u L=180.00n
MM20 net0100 net23 VSS VPW n18 W=0.5u L=180.00n
MM18 net0120 net0100 VSS VPW n18 W=0.5u L=180.00n
MM24 QN net23 VSS VPW n18 W=720.00n L=180.00n
MM6 net0152 c net0139 VNW p18 W=0.58u L=180.00n
MM11 net0132 net0139 VDD VNW p18 W=0.58u L=180.00n
MM12 net0175 net0132 VDD VNW p18 W=0.58u L=180.00n
MM14 net0139 cn net0175 VNW p18 W=580.00n L=180.00n
MM26 net0168 c net23 VNW p18 W=0.49u L=180.00n
MM17 net0132 cn net23 VNW p18 W=0.96u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM5 net0152 D VDD VNW p18 W=0.58u L=180.00n
MM23 net0100 net23 VDD VNW p18 W=1.01u L=180.00n
MM22 net0168 net0100 VDD VNW p18 W=0.73u L=180.00n
MM25 QN net23 VDD VNW p18 W=1.01u L=180.00n
.ENDS DQNUHDV1
.SUBCKT DQNUHDV2 CK D QN VDD VSS VNW VPW
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM12 net127 net180 VDD VNW p18 W=0.59u L=180.00n
MM14 net187 cn net127 VNW p18 W=590.00n L=180.00n
MM26 net120 c net167 VNW p18 W=0.49u L=180.00n
MM17 net180 cn net167 VNW p18 W=0.96u L=180.00n
MM6 net104 c net187 VNW p18 W=0.59u L=180.00n
MM11 net180 net187 VDD VNW p18 W=0.59u L=180.00n
MM5 net104 D VDD VNW p18 W=0.59u L=180.00n
MM23 net148 net167 VDD VNW p18 W=1.01u L=180.00n
MM22 net120 net148 VDD VNW p18 W=0.73u L=180.00n
MM25 QN net167 VDD VNW p18 W=2.02u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM10 net180 net187 VSS VPW n18 W=0.34u L=180.00n
MM13 net187 c net172 VPW n18 W=0.73u L=180.00n
MM15 net172 net180 VSS VPW n18 W=0.34u L=180.00n
MM31 net168 cn net167 VPW n18 W=0.53u L=180.00n
MM20 net148 net167 VSS VPW n18 W=0.53u L=180.00n
MM18 net168 net148 VSS VPW n18 W=0.53u L=180.00n
MM16 net180 c net167 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM4 net152 D VSS VPW n18 W=0.34u L=180.00n
MM24 QN net167 VSS VPW n18 W=1.44u L=180.00n
MM9 net152 cn net187 VPW n18 W=0.51u L=180.00n
.ENDS DQNUHDV2
.SUBCKT DQUHDV0P7 CK D Q VDD VSS VNW VPW
MM24 Q net24 VSS VPW n18 W=0.56u L=180.00n
MM31 net20 cn net15 VPW n18 W=0.5u L=180.00n
MM20 net24 net15 VSS VPW n18 W=0.5u L=180.00n
MM18 net20 net24 VSS VPW n18 W=0.5u L=180.00n
MM16 net40 c net15 VPW n18 W=0.43u L=180.00n
MM15 net32 net40 VSS VPW n18 W=0.36u L=180.00n
MM13 net47 c net32 VPW n18 W=0.73u L=180.00n
MM10 net40 net47 VSS VPW n18 W=0.36u L=180.00n
MM9 net0137 cn net47 VPW n18 W=0.5u L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM4 net0137 D VSS VPW n18 W=0.36u L=180.00n
MM25 Q net24 VDD VNW p18 W=0.79u L=180.00n
MM23 net24 net15 VDD VNW p18 W=1.09u L=180.00n
MM22 net0153 net24 VDD VNW p18 W=0.73u L=180.00n
MM26 net0153 c net15 VNW p18 W=0.49u L=180.00n
MM17 net40 cn net15 VNW p18 W=0.96u L=180.00n
MM14 net47 cn net83 VNW p18 W=580.00n L=180.00n
MM12 net83 net40 VDD VNW p18 W=0.58u L=180.00n
MM11 net40 net47 VDD VNW p18 W=0.58u L=180.00n
MM6 net48 c net47 VNW p18 W=0.58u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM5 net48 D VDD VNW p18 W=0.58u L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
.ENDS DQUHDV0P7
.SUBCKT DQUHDV1 CK D Q VDD VSS VNW VPW
MM9 net0129 cn net55 VPW n18 W=0.5u L=180.00n
MM10 net56 net55 VSS VPW n18 W=0.36u L=180.00n
MM13 net55 c net64 VPW n18 W=0.73u L=180.00n
MM15 net64 net56 VSS VPW n18 W=0.36u L=180.00n
MM31 net0109 cn net79 VPW n18 W=0.5u L=180.00n
MM24 Q net92 VSS VPW n18 W=0.72u L=180.00n
MM16 net56 c net79 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM4 net0129 D VSS VPW n18 W=0.36u L=180.00n
MM20 net92 net79 VSS VPW n18 W=0.5u L=180.00n
MM18 net0109 net92 VSS VPW n18 W=0.5u L=180.00n
MM6 net88 c net55 VNW p18 W=0.58u L=180.00n
MM11 net56 net55 VDD VNW p18 W=0.58u L=180.00n
MM12 net19 net56 VDD VNW p18 W=0.58u L=180.00n
MM14 net55 cn net19 VNW p18 W=580.00n L=180.00n
MM26 net68 c net79 VNW p18 W=0.49u L=180.00n
MM25 Q net92 VDD VNW p18 W=1.01u L=180.00n
MM17 net56 cn net79 VNW p18 W=0.96u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM5 net88 D VDD VNW p18 W=0.58u L=180.00n
MM23 net92 net79 VDD VNW p18 W=1.01u L=180.00n
MM22 net68 net92 VDD VNW p18 W=0.73u L=180.00n
.ENDS DQUHDV1
.SUBCKT DQUHDV2 CK D Q VDD VSS VNW VPW
MM9 net0129 cn net55 VPW n18 W=0.51u L=180.00n
MM10 net56 net55 VSS VPW n18 W=0.34u L=180.00n
MM13 net55 c net64 VPW n18 W=0.73u L=180.00n
MM15 net64 net56 VSS VPW n18 W=0.34u L=180.00n
MM31 net0109 cn net79 VPW n18 W=0.53u L=180.00n
MM24 Q net92 VSS VPW n18 W=1.44u L=180.00n
MM16 net56 c net79 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM4 net0129 D VSS VPW n18 W=0.34u L=180.00n
MM20 net92 net79 VSS VPW n18 W=0.53u L=180.00n
MM18 net0109 net92 VSS VPW n18 W=0.53u L=180.00n
MM6 net88 c net55 VNW p18 W=0.59u L=180.00n
MM11 net56 net55 VDD VNW p18 W=0.59u L=180.00n
MM12 net19 net56 VDD VNW p18 W=0.59u L=180.00n
MM14 net55 cn net19 VNW p18 W=590.00n L=180.00n
MM26 net68 c net79 VNW p18 W=0.49u L=180.00n
MM25 Q net92 VDD VNW p18 W=2.02u L=180.00n
MM17 net56 cn net79 VNW p18 W=0.96u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM5 net88 D VDD VNW p18 W=0.59u L=180.00n
MM23 net92 net79 VDD VNW p18 W=1.01u L=180.00n
MM22 net68 net92 VDD VNW p18 W=0.73u L=180.00n
.ENDS DQUHDV2
.SUBCKT DQUHDV3 CK D Q VDD VSS VNW VPW
MM9 net0129 cn net55 VPW n18 W=0.56u L=180.00n
MM10 net56 net55 VSS VPW n18 W=0.36u L=180.00n
MM13 net55 c net64 VPW n18 W=0.73u L=180.00n
MM15 net64 net56 VSS VPW n18 W=0.36u L=180.00n
MM31 net0109 cn net79 VPW n18 W=0.57u L=180.00n
MM24 Q net92 VSS VPW n18 W=2.16u L=180.00n
MM16 net56 c net79 VPW n18 W=0.43u L=180.00n
MM0 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 c cn VSS VPW n18 W=250.00n L=180.00n
MM4 net0129 D VSS VPW n18 W=0.36u L=180.00n
MM20 net92 net79 VSS VPW n18 W=0.57u L=180.00n
MM18 net0109 net92 VSS VPW n18 W=0.57u L=180.00n
MM6 net88 c net55 VNW p18 W=0.58u L=180.00n
MM11 net56 net55 VDD VNW p18 W=0.51u L=180.00n
MM12 net19 net56 VDD VNW p18 W=0.51u L=180.00n
MM14 net55 cn net19 VNW p18 W=0.51u L=180.00n
MM26 net68 c net79 VNW p18 W=0.49u L=180.00n
MM25 Q net92 VDD VNW p18 W=3.03u L=180.00n
MM17 net56 cn net79 VNW p18 W=0.49u L=180.00n
MM1 cn CK VDD VNW p18 W=250.00n L=180.00n
MM3 c cn VDD VNW p18 W=420.00n L=180.00n
MM5 net88 D VDD VNW p18 W=0.58u L=180.00n
MM23 net92 net79 VDD VNW p18 W=1.01u L=180.00n
MM22 net68 net92 VDD VNW p18 W=0.66u L=180.00n
.ENDS DQUHDV3
.SUBCKT DRNQUHDV0P7 CK D Q RDN VDD VSS VNW VPW
MM27 net_0167 net4 VSS VPW n18 W=0.42u L=180.00n
MM25 net8 c net9 VPW n18 W=0.715u L=180.00n
MM23 net9 RDN net_97 VPW n18 W=0.28u L=180.00n
MM22 net_97 net12 VSS VPW n18 W=0.28u L=180.00n
MM15 net12 c net11 VPW n18 W=0.42u L=180.00n
MM12 net12 net8 VSS VPW n18 W=280.00n L=180.00n
MM9 net7 cn net8 VPW n18 W=0.43u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM3 cn CK VSS VPW n18 W=420.00n L=180.00n
MM1 net7 D VSS VPW n18 W=0.37u L=180.00n
MM11 net11 cn net_0167 VPW n18 W=0.42u L=180.00n
MM19 net4 net11 net_81 VPW n18 W=0.42u L=180.00n
MM18 net_81 RDN VSS VPW n18 W=0.42u L=180.00n
MM4 Q net4 VSS VPW n18 W=0.56u L=180.00n
MM26 net14 net4 VDD VNW p18 W=0.28u L=180.00n
MM24 net8 cn net_0195 VNW p18 W=0.495u L=180.00n
MM21 net_0195 net12 VDD VNW p18 W=0.335u L=180.00n
MM20 net_0195 RDN VDD VNW p18 W=0.46u L=180.00n
MM14 net12 cn net11 VNW p18 W=430.00n L=180.00n
MM10 net12 net8 VDD VNW p18 W=0.37u L=180.00n
MM8 net_0220 c net8 VNW p18 W=0.495u L=180.00n
MM6 c cn VDD VNW p18 W=0.42u L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM13 net11 c net14 VNW p18 W=0.28u L=180.00n
MM0 net_0220 D VDD VNW p18 W=0.495u L=180.00n
MM16 net4 RDN VDD VNW p18 W=1.045u L=180.00n
MM17 net4 net11 VDD VNW p18 W=1.09u L=180.00n
MM5 Q net4 VDD VNW p18 W=0.81u L=180.00n
.ENDS DRNQUHDV0P7
.SUBCKT DRNQUHDV1 CK D Q RDN VDD VSS VNW VPW
MM1 net7 D VSS VPW n18 W=0.28u L=180.00n
MM9 net7 cn net8 VPW n18 W=0.28u L=180.00n
MM12 net12 net8 VSS VPW n18 W=0.28u L=180.00n
MM15 net12 c net11 VPW n18 W=0.42u L=180.00n
MM22 net_21 net12 VSS VPW n18 W=0.25u L=180.00n
MM23 net_0148 RDN net_21 VPW n18 W=0.25u L=180.00n
MM25 net8 c net_0148 VPW n18 W=0.25u L=180.00n
MM19 net4 net11 net_37 VPW n18 W=0.42u L=180.00n
MM18 net_37 RDN VSS VPW n18 W=0.42u L=180.00n
MM4 Q net4 VSS VPW n18 W=0.72u L=180.00n
MM27 net_0169 net4 VSS VPW n18 W=0.42u L=180.00n
MM11 net11 cn net_0169 VPW n18 W=0.42u L=180.00n
MM3 cn CK VSS VPW n18 W=0.42u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM0 net_0178 D VDD VNW p18 W=0.495u L=180.00n
MM8 net_0178 c net8 VNW p18 W=0.495u L=180.00n
MM10 net12 net8 VDD VNW p18 W=0.37u L=180.00n
MM14 net12 cn net11 VNW p18 W=0.43u L=180.00n
MM20 net9 RDN VDD VNW p18 W=0.42u L=180.00n
MM21 net9 net12 VDD VNW p18 W=0.335u L=180.00n
MM24 net8 cn net9 VNW p18 W=0.42u L=180.00n
MM17 net4 net11 VDD VNW p18 W=1.01u L=180.00n
MM16 net4 RDN VDD VNW p18 W=1.01u L=180.00n
MM5 Q net4 VDD VNW p18 W=1.01u L=180.00n
MM26 net14 net4 VDD VNW p18 W=0.28u L=180.00n
MM13 net11 c net14 VNW p18 W=0.28u L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM6 c cn VDD VNW p18 W=0.42u L=180.00n
.ENDS DRNQUHDV1
.SUBCKT DRNQUHDV2 CK D Q RDN VDD VSS VNW VPW
MM1 net_0124 D VSS VPW n18 W=0.28u L=180.00n
MM9 net_0124 cn net8 VPW n18 W=0.28u L=180.00n
MM12 net12 net8 VSS VPW n18 W=0.28u L=180.00n
MM15 net12 c net11 VPW n18 W=0.42u L=180.00n
MM22 net_21 net12 VSS VPW n18 W=0.25u L=180.00n
MM23 net_0151 RDN net_21 VPW n18 W=0.25u L=180.00n
MM25 net8 c net_0151 VPW n18 W=0.25u L=180.00n
MM19 net4 net11 net_37 VPW n18 W=0.42u L=180.00n
MM18 net_37 RDN VSS VPW n18 W=0.42u L=180.00n
MM4 Q net4 VSS VPW n18 W=1.44u L=180.00n
MM27 net14 net4 VSS VPW n18 W=0.42u L=180.00n
MM11 net11 cn net14 VPW n18 W=0.42u L=180.00n
MM3 cn CK VSS VPW n18 W=0.42u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM0 net7 D VDD VNW p18 W=0.495u L=180.00n
MM8 net7 c net8 VNW p18 W=0.495u L=180.00n
MM10 net12 net8 VDD VNW p18 W=0.37u L=180.00n
MM14 net12 cn net11 VNW p18 W=0.43u L=180.00n
MM20 net9 RDN VDD VNW p18 W=0.42u L=180.00n
MM21 net9 net12 VDD VNW p18 W=0.335u L=180.00n
MM24 net8 cn net9 VNW p18 W=0.42u L=180.00n
MM17 net4 net11 VDD VNW p18 W=1.01u L=180.00n
MM16 net4 RDN VDD VNW p18 W=1.01u L=180.00n
MM5 Q net4 VDD VNW p18 W=2.02u L=180.00n
MM26 net_0227 net4 VDD VNW p18 W=0.28u L=180.00n
MM13 net11 c net_0227 VNW p18 W=0.28u L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM6 c cn VDD VNW p18 W=0.42u L=180.00n
.ENDS DRNQUHDV2
.SUBCKT DRNQUHDV3 CK D Q RDN VDD VSS VNW VPW
MM1 net7 D VSS VPW n18 W=0.28u L=180.00n
MM9 net7 cn net8 VPW n18 W=0.28u L=180.00n
MM12 net12 net8 VSS VPW n18 W=0.28u L=180.00n
MM15 net12 c net11 VPW n18 W=0.42u L=180.00n
MM22 net_21 net12 VSS VPW n18 W=0.25u L=180.00n
MM23 net9 RDN net_21 VPW n18 W=0.25u L=180.00n
MM25 net8 c net9 VPW n18 W=0.25u L=180.00n
MM19 net4 net11 net_37 VPW n18 W=0.42u L=180.00n
MM18 net_37 RDN VSS VPW n18 W=0.42u L=180.00n
MM4 Q net4 VSS VPW n18 W=2.16u L=180.00n
MM27 net14 net4 VSS VPW n18 W=0.42u L=180.00n
MM11 net11 cn net14 VPW n18 W=0.42u L=180.00n
MM3 cn CK VSS VPW n18 W=0.42u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM0 net_0180 D VDD VNW p18 W=0.495u L=180.00n
MM8 net_0180 c net8 VNW p18 W=0.495u L=180.00n
MM10 net12 net8 VDD VNW p18 W=0.37u L=180.00n
MM14 net12 cn net11 VNW p18 W=0.43u L=180.00n
MM20 net_0207 RDN VDD VNW p18 W=0.42u L=180.00n
MM21 net_0207 net12 VDD VNW p18 W=0.335u L=180.00n
MM24 net8 cn net_0207 VNW p18 W=0.42u L=180.00n
MM17 net4 net11 VDD VNW p18 W=1.01u L=180.00n
MM16 net4 RDN VDD VNW p18 W=1.01u L=180.00n
MM5 Q net4 VDD VNW p18 W=3.03u L=180.00n
MM26 net_0227 net4 VDD VNW p18 W=0.28u L=180.00n
MM13 net11 c net_0227 VNW p18 W=0.28u L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM6 c cn VDD VNW p18 W=0.42u L=180.00n
.ENDS DRNQUHDV3
****Sub-Circuit for DRQUHDV0P7, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT DRQUHDV0P7 CK D Q RD VDD VSS VNW VPW
MM22 Q net47 VSS VPW n18 W=560.00n L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM0 net17 cn net13 VPW n18 W=420.00n L=180.00n
MM1 net13 D VSS VPW n18 W=420.00n L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=420.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 net84 D VDD VNW p18 W=560.00n L=180.00n
MM3 net17 c net84 VNW p18 W=560.00n L=180.00n
MM23 Q net47 VDD VNW p18 W=790.00n L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=790.00n L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
.ENDS DRQUHDV0P7
****Sub-Circuit for DRQUHDV1, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT DRQUHDV1 CK D Q RD VDD VSS VNW VPW
MM22 Q net47 VSS VPW n18 W=720.00n L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM0 net17 cn net13 VPW n18 W=420.00n L=180.00n
MM1 net13 D VSS VPW n18 W=420.00n L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=560.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 net84 D VDD VNW p18 W=560.00n L=180.00n
MM3 net17 c net84 VNW p18 W=560.00n L=180.00n
MM23 Q net47 VDD VNW p18 W=1.01u L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=1.01u L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
.ENDS DRQUHDV1
****Sub-Circuit for DRQUHDV2, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT DRQUHDV2 CK D Q RD VDD VSS VNW VPW
MM22 Q net47 VSS VPW n18 W=1.44u L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM0 net17 cn net13 VPW n18 W=420.00n L=180.00n
MM1 net13 D VSS VPW n18 W=420.00n L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=560.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 net84 D VDD VNW p18 W=560.00n L=180.00n
MM3 net17 c net84 VNW p18 W=560.00n L=180.00n
MM23 Q net47 VDD VNW p18 W=2.02u L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=1.01u L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
.ENDS DRQUHDV2
****Sub-Circuit for DRQUHDV3, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT DRQUHDV3 CK D Q RD VDD VSS VNW VPW
MM22 Q net47 VSS VPW n18 W=2.16u L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM0 net17 cn net13 VPW n18 W=420.00n L=180.00n
MM1 net13 D VSS VPW n18 W=420.00n L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=560.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM2 net84 D VDD VNW p18 W=560.00n L=180.00n
MM3 net17 c net84 VNW p18 W=560.00n L=180.00n
MM23 Q net47 VDD VNW p18 W=3.03u L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=1.01u L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
.ENDS DRQUHDV3
.SUBCKT DSNQUHDV0P7 CK D Q SDN VDD VSS VNW VPW
MM20 net7 D VSS VPW n18 W=0.63u L=180.00n
MM22 cn CK VSS VPW n18 W=420.00n L=180.00n
MM14 net_0134 net10 VSS VPW n18 W=0.43u L=180.00n
MM11 net7 cn net6 VPW n18 W=0.48u L=180.00n
MM10 net_0134 c net6 VPW n18 W=0.4u L=180.00n
MM4 Q net4 VSS VPW n18 W=0.56u L=180.00n
MM19 net10 net6 net_41 VPW n18 W=0.4u L=180.00n
MM18 net_41 SDN VSS VPW n18 W=0.4u L=180.00n
MM0 net4 net12 VSS VPW n18 W=0.51u L=180.00n
MM9 net11 SDN net_49 VPW n18 W=0.4u L=180.00n
MM8 net_49 net4 VSS VPW n18 W=0.4u L=180.00n
MM6 c cn VSS VPW n18 W=420.00n L=180.00n
MM38 net10 c net12 VPW n18 W=0.4u L=180.00n
MM37 net11 cn net12 VPW n18 W=0.4u L=180.00n
MM23 cn CK VDD VNW p18 W=250.00n L=180.00n
MM21 net7 D VDD VNW p18 W=1.01u L=180.00n
MM15 net8 net10 VDD VNW p18 W=0.435u L=180.00n
MM13 net7 c net6 VNW p18 W=0.435u L=180.00n
MM12 net8 cn net6 VNW p18 W=435.00n L=180.00n
MM5 Q net4 VDD VNW p18 W=0.79u L=180.00n
MM17 net10 net6 VDD VNW p18 W=0.495u L=180.00n
MM16 net10 SDN VDD VNW p18 W=0.495u L=180.00n
MM1 net4 net12 VDD VNW p18 W=1.01u L=180.00n
MM3 net11 net4 VDD VNW p18 W=0.755u L=180.00n
MM2 net11 SDN VDD VNW p18 W=0.96u L=180.00n
MM7 c cn VDD VNW p18 W=420.00n L=180.00n
MM39 net10 cn net12 VNW p18 W=0.73u L=180.00n
MM40 net11 c net12 VNW p18 W=0.72u L=180.00n
.ENDS DSNQUHDV0P7
.SUBCKT DSNQUHDV1 CK D Q SDN VDD VSS VNW VPW
MM9 net11 SDN net_227 VPW n18 W=0.4u L=180.00n
MM8 net_227 net4 VSS VPW n18 W=0.4u L=180.00n
MM37 net11 cn net12 VPW n18 W=0.4u L=180.00n
MM4 Q net4 VSS VPW n18 W=0.72u L=180.00n
MM0 net4 net12 VSS VPW n18 W=0.51u L=180.00n
MM38 net10 c net12 VPW n18 W=0.4u L=180.00n
MM19 net10 net6 net_203 VPW n18 W=0.4u L=180.00n
MM18 net_203 SDN VSS VPW n18 W=0.4u L=180.00n
MM22 cn CK VSS VPW n18 W=420.00n L=180.00n
MM6 c cn VSS VPW n18 W=420.00n L=180.00n
MM14 net_0170 net10 VSS VPW n18 W=0.43u L=180.00n
MM20 net_0222 D VSS VPW n18 W=0.6u L=180.00n
MM11 net_0222 cn net6 VPW n18 W=0.48u L=180.00n
MM10 net_0170 c net6 VPW n18 W=0.4u L=180.00n
MM3 net11 net4 VDD VNW p18 W=0.755u L=180.00n
MM2 net11 SDN VDD VNW p18 W=0.96u L=180.00n
MM40 net11 c net12 VNW p18 W=0.72u L=180.00n
MM5 Q net4 VDD VNW p18 W=1.01u L=180.00n
MM1 net4 net12 VDD VNW p18 W=1.01u L=180.00n
MM39 net10 cn net12 VNW p18 W=0.73u L=180.00n
MM17 net10 net6 VDD VNW p18 W=0.495u L=180.00n
MM16 net10 SDN VDD VNW p18 W=0.495u L=180.00n
MM23 cn CK VDD VNW p18 W=250.00n L=180.00n
MM7 c cn VDD VNW p18 W=420.00n L=180.00n
MM15 net8 net10 VDD VNW p18 W=0.435u L=180.00n
MM12 net8 cn net6 VNW p18 W=435.00n L=180.00n
MM21 net_0222 D VDD VNW p18 W=1.01u L=180.00n
MM13 net_0222 c net6 VNW p18 W=0.435u L=180.00n
.ENDS DSNQUHDV1
.SUBCKT DSNQUHDV2 CK D Q SDN VDD VSS VNW VPW
MM4 Q net4 VSS VPW n18 W=1.44u L=180.00n
MM0 net4 net12 VSS VPW n18 W=0.51u L=180.00n
MM38 net10 c net12 VPW n18 W=0.4u L=180.00n
MM19 net10 net6 net_203 VPW n18 W=0.4u L=180.00n
MM18 net_203 SDN VSS VPW n18 W=0.4u L=180.00n
MM22 cn CK VSS VPW n18 W=420.00n L=180.00n
MM6 c cn VSS VPW n18 W=420.00n L=180.00n
MM14 net_0150 net10 VSS VPW n18 W=0.43u L=180.00n
MM10 net_0150 c net6 VPW n18 W=0.4u L=180.00n
MM20 net_0154 D VSS VPW n18 W=0.6u L=180.00n
MM11 net_0154 cn net6 VPW n18 W=0.48u L=180.00n
MM9 net11 SDN net_227 VPW n18 W=0.4u L=180.00n
MM8 net_227 net4 VSS VPW n18 W=0.4u L=180.00n
MM37 net11 cn net12 VPW n18 W=0.4u L=180.00n
MM3 net11 net4 VDD VNW p18 W=0.755u L=180.00n
MM2 net11 SDN VDD VNW p18 W=0.96u L=180.00n
MM40 net11 c net12 VNW p18 W=0.72u L=180.00n
MM5 Q net4 VDD VNW p18 W=2.02u L=180.00n
MM1 net4 net12 VDD VNW p18 W=1.01u L=180.00n
MM39 net10 cn net12 VNW p18 W=0.73u L=180.00n
MM17 net10 net6 VDD VNW p18 W=0.495u L=180.00n
MM16 net10 SDN VDD VNW p18 W=0.495u L=180.00n
MM23 cn CK VDD VNW p18 W=250.00n L=180.00n
MM7 c cn VDD VNW p18 W=420.00n L=180.00n
MM15 net8 net10 VDD VNW p18 W=0.435u L=180.00n
MM12 net8 cn net6 VNW p18 W=435.00n L=180.00n
MM21 net_0154 D VDD VNW p18 W=1.01u L=180.00n
MM13 net_0154 c net6 VNW p18 W=0.435u L=180.00n
.ENDS DSNQUHDV2
.SUBCKT DSNQUHDV3 CK D Q SDN VDD VSS VNW VPW
MM4 Q net4 VSS VPW n18 W=2.16u L=180.00n
MM0 net4 net12 VSS VPW n18 W=0.51u L=180.00n
MM38 net10 c net12 VPW n18 W=0.4u L=180.00n
MM19 net10 net6 net_203 VPW n18 W=0.4u L=180.00n
MM18 net_203 SDN VSS VPW n18 W=0.4u L=180.00n
MM22 cn CK VSS VPW n18 W=420.00n L=180.00n
MM6 c cn VSS VPW n18 W=420.00n L=180.00n
MM14 net8 net10 VSS VPW n18 W=0.43u L=180.00n
MM10 net8 c net6 VPW n18 W=0.4u L=180.00n
MM20 net_0222 D VSS VPW n18 W=0.6u L=180.00n
MM11 net_0222 cn net6 VPW n18 W=0.48u L=180.00n
MM9 net11 SDN net_227 VPW n18 W=0.4u L=180.00n
MM8 net_227 net4 VSS VPW n18 W=0.4u L=180.00n
MM37 net11 cn net12 VPW n18 W=0.4u L=180.00n
MM3 net11 net4 VDD VNW p18 W=0.755u L=180.00n
MM2 net11 SDN VDD VNW p18 W=0.96u L=180.00n
MM40 net11 c net12 VNW p18 W=0.72u L=180.00n
MM5 Q net4 VDD VNW p18 W=3.03u L=180.00n
MM1 net4 net12 VDD VNW p18 W=1.01u L=180.00n
MM39 net10 cn net12 VNW p18 W=0.73u L=180.00n
MM17 net10 net6 VDD VNW p18 W=0.495u L=180.00n
MM16 net10 SDN VDD VNW p18 W=0.495u L=180.00n
MM23 cn CK VDD VNW p18 W=250.00n L=180.00n
MM7 c cn VDD VNW p18 W=420.00n L=180.00n
MM15 net_0218 net10 VDD VNW p18 W=0.435u L=180.00n
MM12 net_0218 cn net6 VNW p18 W=435.00n L=180.00n
MM21 net_0222 D VDD VNW p18 W=1.01u L=180.00n
MM13 net_0222 c net6 VNW p18 W=0.435u L=180.00n
.ENDS DSNQUHDV3
.SUBCKT DSRNQUHDV1 CK D Q RDN SDN VDD VSS VNW VPW
MM28 net81 cn net129 VPW n18 W=0.445u L=180.00n
MM39 net77 net113 VSS VPW n18 W=0.42u L=180.00n
MM38 net73 SDN net77 VPW n18 W=0.42u L=180.00n
MM33 net81 c net105 VPW n18 W=0.445u L=180.00n
MM31 net121 net81 VSS VPW n18 W=0.49u L=180.00n
MM19 net113 net100 net117 VPW n18 W=0.53u L=180.00n
MM23 net105 RDN net125 VPW n18 W=0.445u L=180.00n
MM37 net100 cn net73 VPW n18 W=0.42u L=180.00n
MM15 net93 c net100 VPW n18 W=0.42u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM3 cn CK VSS VPW n18 W=420.00n L=180.00n
MM12 net93 SDN net121 VPW n18 W=0.49u L=180.00n
MM18 net117 RDN VSS VPW n18 W=0.53u L=180.00n
MM4 Q net113 VSS VPW n18 W=0.72u L=180.00n
MM1 net129 D VSS VPW n18 W=0.445u L=180.00n
MM22 net125 net93 VSS VPW n18 W=0.445u L=180.00n
MM29 net81 c net136 VNW p18 W=0.42u L=180.00n
MM34 net137 net113 VDD VNW p18 W=0.42u L=180.00n
MM5 Q net113 VDD VNW p18 W=1.01u L=180.00n
MM17 net113 net100 VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net137 VNW p18 W=0.425u L=180.00n
MM16 net113 RDN VDD VNW p18 W=0.42u L=180.00n
MM0 net136 D VDD VNW p18 W=0.42u L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM6 c cn VDD VNW p18 W=0.42u L=180.00n
MM10 net93 net81 VDD VNW p18 W=0.42u L=180.00n
MM14 net93 cn net100 VNW p18 W=0.425u L=180.00n
MM20 net153 RDN VDD VNW p18 W=0.42u L=180.00n
MM21 net153 net93 VDD VNW p18 W=0.42u L=180.00n
MM32 net81 cn net153 VNW p18 W=0.42u L=180.00n
MM30 net93 SDN VDD VNW p18 W=0.37u L=180.00n
MM35 net137 SDN VDD VNW p18 W=0.42u L=180.00n
.ENDS DSRNQUHDV1
.SUBCKT DSRNQUHDV2 CK D Q RDN SDN VDD VSS VNW VPW
MM28 net81 cn net129 VPW n18 W=0.445u L=180.00n
MM39 net77 net113 VSS VPW n18 W=0.42u L=180.00n
MM38 net73 SDN net77 VPW n18 W=0.42u L=180.00n
MM33 net81 c net105 VPW n18 W=0.445u L=180.00n
MM1 net129 D VSS VPW n18 W=0.445u L=180.00n
MM22 net125 net93 VSS VPW n18 W=0.445u L=180.00n
MM31 net121 net81 VSS VPW n18 W=0.49u L=180.00n
MM18 net117 RDN VSS VPW n18 W=0.53u L=180.00n
MM19 net113 net100 net117 VPW n18 W=0.53u L=180.00n
MM37 net100 cn net73 VPW n18 W=0.42u L=180.00n
MM23 net105 RDN net125 VPW n18 W=0.445u L=180.00n
MM4 Q net113 VSS VPW n18 W=1.44u L=180.00n
MM15 net93 c net100 VPW n18 W=0.42u L=180.00n
MM12 net93 SDN net121 VPW n18 W=0.49u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM3 cn CK VSS VPW n18 W=420.00n L=180.00n
MM30 net93 SDN VDD VNW p18 W=0.37u L=180.00n
MM35 net137 SDN VDD VNW p18 W=0.42u L=180.00n
MM34 net137 net113 VDD VNW p18 W=0.42u L=180.00n
MM29 net81 c net136 VNW p18 W=0.42u L=180.00n
MM5 Q net113 VDD VNW p18 W=2.02u L=180.00n
MM17 net113 net100 VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net137 VNW p18 W=0.425u L=180.00n
MM16 net113 RDN VDD VNW p18 W=0.42u L=180.00n
MM0 net136 D VDD VNW p18 W=0.42u L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM6 c cn VDD VNW p18 W=0.42u L=180.00n
MM10 net93 net81 VDD VNW p18 W=0.42u L=180.00n
MM14 net93 cn net100 VNW p18 W=0.425u L=180.00n
MM20 net153 RDN VDD VNW p18 W=0.42u L=180.00n
MM21 net153 net93 VDD VNW p18 W=0.42u L=180.00n
MM32 net81 cn net153 VNW p18 W=0.42u L=180.00n
.ENDS DSRNQUHDV2
.SUBCKT FDCAPUHD12 VDD VSS VNW VPW
MM36 net1 net3 VSS VPW n18 W=720.00n L=5.33u
MM31 net3 net1 VDD VNW p18 W=1.01u L=5.33u
.ENDS FDCAPUHD12
.SUBCKT FDCAPUHD16 VDD VSS VNW VPW
MM36 net1 net3 VSS VPW n18 W=720.00n L=7.57u
MM31 net3 net1 VDD VNW p18 W=1.01u L=7.57u
.ENDS FDCAPUHD16
.SUBCKT FDCAPUHD24 VDD VSS VNW VPW
MM36 net1 net3 VSS VPW n18 W=720.00n L=12.05u
MM31 net3 net1 VDD VNW p18 W=1.01u L=12.05u
.ENDS FDCAPUHD24
.SUBCKT FDCAPUHD32 VDD VSS VNW VPW
MM36 net1 net3 VSS VPW n18 W=720.00n L=16.53u
MM31 net3 net1 VDD VNW p18 W=1.01u L=16.53u
.ENDS FDCAPUHD32
.SUBCKT FDCAPUHD4 VDD VSS VNW VPW
MM36 net1 net3 VSS VPW n18 W=660.00n L=1000.00n
MM31 net3 net1 VDD VNW p18 W=1.01u L=1000.00n
.ENDS FDCAPUHD4
.SUBCKT FDCAPUHD64 VDD VSS VNW VPW
MM36 net1 net3 VSS VPW n18 W=720.00n L=34.45u
MM31 net3 net1 VDD VNW p18 W=1.01u L=34.45u
.ENDS FDCAPUHD64
.SUBCKT FDCAPUHD8 VDD VSS VNW VPW
MM31 net7 net5 VDD VNW p18 W=1.01u L=3.09u
MM36 net5 net7 VSS VPW n18 W=720.00n L=3.09u
.ENDS FDCAPUHD8
.SUBCKT FILLTIEUHD VDD VSS
.ENDS FILLTIEUHD
.SUBCKT F_DIODENUHD2 A VDD VSS VNW VPW
DD1 VPW A ndio18 AREA=0.672p PJ=3.28u
.ENDS F_DIODENUHD2
.SUBCKT F_DIODEUHD2 A VDD VSS VNW VPW
DD0 A VNW pdio18 AREA=0.8484p PJ=3.7u
DD1 VPW A ndio18 AREA=0.672p PJ=3.28u
.ENDS F_DIODEUHD2
.SUBCKT F_FILLUHD1 VDD VSS VNW VPW
.ENDS F_FILLUHD1
.SUBCKT F_FILLUHD16 VDD VSS VNW VPW
.ENDS F_FILLUHD16
.SUBCKT F_FILLUHD2 VDD VSS VNW VPW
.ENDS F_FILLUHD2
.SUBCKT F_FILLUHD32 VDD VSS VNW VPW
.ENDS F_FILLUHD32
.SUBCKT F_FILLUHD4 VDD VSS VNW VPW
.ENDS F_FILLUHD4
.SUBCKT F_FILLUHD8 VDD VSS VNW VPW
.ENDS F_FILLUHD8
.SUBCKT INUHDV0P4 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=0.28u L=180.00n
MM13 ZN I VDD VNW p18 W=490.0n L=180.00n
.ENDS INUHDV0P4
.SUBCKT INUHDV0P7 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=560.00n L=180.00n
MM13 ZN I VDD VNW p18 W=790.0n L=180.00n
.ENDS INUHDV0P7
.SUBCKT INUHDV1 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=720.00n L=180.00n
MM13 ZN I VDD VNW p18 W=1.01u L=180.00n
.ENDS INUHDV1
.SUBCKT INUHDV16 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=11.52u L=180.00n
MM13 ZN I VDD VNW p18 W=16.16u L=180.00n
.ENDS INUHDV16
.SUBCKT INUHDV2 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=1.44u L=180.00n
MM13 ZN I VDD VNW p18 W=2.02u L=180.00n
.ENDS INUHDV2
.SUBCKT INUHDV20 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=14.4u L=180.00n
MM13 ZN I VDD VNW p18 W=20.2u L=180.00n
.ENDS INUHDV20
.SUBCKT INUHDV24 I ZN VDD VSS VNW VPW
MM13 ZN I VDD VNW p18 W=24.24u L=180.00n
MM12 ZN I VSS VPW n18 W=17.28u L=180.00n
.ENDS INUHDV24
.SUBCKT INUHDV3 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=2.16u L=180.00n
MM13 ZN I VDD VNW p18 W=3.03u L=180.00n
.ENDS INUHDV3
.SUBCKT INUHDV4 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=2.88u L=180.00n
MM13 ZN I VDD VNW p18 W=4.04u L=180.00n
.ENDS INUHDV4
.SUBCKT INUHDV6 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=4.32u L=180.00n
MM13 ZN I VDD VNW p18 W=6.06u L=180.00n
.ENDS INUHDV6
.SUBCKT INUHDV8 I ZN VDD VSS VNW VPW
MM12 ZN I VSS VPW n18 W=5.76u L=180.00n
MM13 ZN I VDD VNW p18 W=8.08u L=180.00n
.ENDS INUHDV8
.SUBCKT LAHQUHDV0P7 D E Q VDD VSS VNW VPW
MM9 c E VSS VPW n18 W=430.00n L=180.00n
MM6 cn c VSS VPW n18 W=720.00n L=180.00n
MM4 net24 net28 VSS VPW n18 W=0.435u L=180.00n
MM0 net32 D VSS VPW n18 W=0.42u L=180.00n
MM1 net28 cn net32 VPW n18 W=0.42u L=180.00n
MM25 Q net28 VSS VPW n18 W=0.565u L=180.00n
MM22 net16 net24 VSS VPW n18 W=0.42u L=180.00n
MM23 net28 c net16 VPW n18 W=0.42u L=180.00n
MM8 c E VDD VNW p18 W=0.59u L=180.00n
MM7 cn c VDD VNW p18 W=0.95u L=180.00n
MM5 net24 net28 VDD VNW p18 W=0.59u L=180.00n
MM3 net67 D VDD VNW p18 W=0.575u L=180.00n
MM2 net28 c net67 VNW p18 W=0.59u L=180.00n
MM24 Q net28 VDD VNW p18 W=0.795u L=180.00n
MM20 net28 cn net51 VNW p18 W=0.585u L=180.00n
MM21 net51 net24 VDD VNW p18 W=0.585u L=180.00n
.ENDS LAHQUHDV0P7
.SUBCKT LAHQUHDV1 D E Q VDD VSS VNW VPW
MM2 net40 c net7 VNW p18 W=0.59u L=180.00n
MM3 net7 D VDD VNW p18 W=0.59u L=180.00n
MM5 net44 net40 VDD VNW p18 W=0.585u L=180.00n
MM21 net23 net44 VDD VNW p18 W=0.59u L=180.00n
MM20 net40 cn net23 VNW p18 W=0.59u L=180.00n
MM24 Q net40 VDD VNW p18 W=1.01u L=180.00n
MM7 cn c VDD VNW p18 W=1.01u L=180.00n
MM8 c E VDD VNW p18 W=0.59u L=180.00n
MM0 net36 D VSS VPW n18 W=430.00n L=180.00n
MM1 net40 cn net36 VPW n18 W=430.00n L=180.00n
MM4 net44 net40 VSS VPW n18 W=0.44u L=180.00n
MM23 net40 c net52 VPW n18 W=430.00n L=180.00n
MM22 net52 net44 VSS VPW n18 W=430.00n L=180.00n
MM25 Q net40 VSS VPW n18 W=720.00n L=180.00n
MM6 cn c VSS VPW n18 W=0.67u L=180.00n
MM9 c E VSS VPW n18 W=430.00n L=180.00n
.ENDS LAHQUHDV1
.SUBCKT LAHQUHDV2 D E Q VDD VSS VNW VPW
MM2 net40 c net7 VNW p18 W=0.945u L=180.00n
MM3 net7 D VDD VNW p18 W=0.945u L=180.00n
MM5 net44 net40 VDD VNW p18 W=0.585u L=180.00n
MM21 net23 net44 VDD VNW p18 W=0.585u L=180.00n
MM20 net40 cn net23 VNW p18 W=0.585u L=180.00n
MM24 Q net40 VDD VNW p18 W=2.02u L=180.00n
MM7 cn c VDD VNW p18 W=1.01u L=180.00n
MM8 c E VDD VNW p18 W=0.59u L=180.00n
MM0 net36 D VSS VPW n18 W=0.635u L=180.00n
MM1 net40 cn net36 VPW n18 W=0.635u L=180.00n
MM4 net44 net40 VSS VPW n18 W=0.435u L=180.00n
MM23 net40 c net52 VPW n18 W=0.435u L=180.00n
MM22 net52 net44 VSS VPW n18 W=0.435u L=180.00n
MM25 Q net40 VSS VPW n18 W=1.44u L=180.00n
MM6 cn c VSS VPW n18 W=0.67u L=180.00n
MM9 c E VSS VPW n18 W=430.00n L=180.00n
.ENDS LAHQUHDV2
.SUBCKT LAHQUHDV3 D E Q VDD VSS VNW VPW
MM9 c E VSS VPW n18 W=430.00n L=180.00n
MM6 cn c VSS VPW n18 W=0.67u L=180.00n
MM25 Q net28 VSS VPW n18 W=2.16u L=180.00n
MM22 net16 net24 VSS VPW n18 W=0.435u L=180.00n
MM23 net28 c net16 VPW n18 W=0.435u L=180.00n
MM4 net24 net28 VSS VPW n18 W=0.435u L=180.00n
MM1 net28 cn net32 VPW n18 W=0.635u L=180.00n
MM0 net32 D VSS VPW n18 W=0.635u L=180.00n
MM8 c E VDD VNW p18 W=0.59u L=180.00n
MM7 cn c VDD VNW p18 W=1.01u L=180.00n
MM24 Q net28 VDD VNW p18 W=3.03u L=180.00n
MM20 net28 cn net51 VNW p18 W=0.585u L=180.00n
MM21 net51 net24 VDD VNW p18 W=0.585u L=180.00n
MM5 net24 net28 VDD VNW p18 W=0.585u L=180.00n
MM3 net67 D VDD VNW p18 W=0.945u L=180.00n
MM2 net28 c net67 VNW p18 W=0.945u L=180.00n
.ENDS LAHQUHDV3
.SUBCKT LAHRNQUHDV0P7 D E Q RDN VDD VSS VNW VPW
MM6 en E VSS VPW n18 W=430.00n L=180.00n
MM4 enn en VSS VPW n18 W=430.00n L=180.00n
MM18 net_13 RDN VSS VPW n18 W=0.43u L=180.00n
MM17 net_17 D net_13 VPW n18 W=0.43u L=180.00n
MM15 net_21 net5 net_25 VPW n18 W=0.42u L=180.00n
MM14 net_25 RDN VSS VPW n18 W=0.42u L=180.00n
MM19 net_69 enn net_17 VPW n18 W=0.43u L=180.00n
MM20 net_69 en net_21 VPW n18 W=0.42u L=180.00n
MM2 net5 net_69 VSS VPW n18 W=0.435u L=180.00n
MM0 Q net_69 VSS VPW n18 W=560.00n L=180.00n
MM7 en E VDD VNW p18 W=0.96u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM8 net_69 RDN VDD VNW p18 W=0.505u L=180.00n
MM13 net_64 net5 VDD VNW p18 W=0.95u L=180.00n
MM11 net_69 enn net_64 VNW p18 W=0.95u L=180.00n
MM10 net_72 D VDD VNW p18 W=0.52u L=180.00n
MM9 net_69 en net_72 VNW p18 W=0.76u L=180.00n
MM3 net5 net_69 VDD VNW p18 W=490.0n L=180.00n
MM1 Q net_69 VDD VNW p18 W=0.8u L=180.00n
.ENDS LAHRNQUHDV0P7
.SUBCKT LAHRNQUHDV1 D E Q RDN VDD VSS VNW VPW
MM1 Q net7 VDD VNW p18 W=1.01u L=180.00n
MM3 net5 net7 VDD VNW p18 W=490.0n L=180.00n
MM8 net7 RDN VDD VNW p18 W=0.505u L=180.00n
MM9 net7 en net_16 VNW p18 W=0.76u L=180.00n
MM10 net_16 D VDD VNW p18 W=0.52u L=180.00n
MM11 net7 enn net_20 VNW p18 W=0.95u L=180.00n
MM13 net_20 net5 VDD VNW p18 W=0.95u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM7 en E VDD VNW p18 W=0.96u L=180.00n
MM20 net7 en net_61 VPW n18 W=0.42u L=180.00n
MM19 net7 enn net_45 VPW n18 W=0.43u L=180.00n
MM0 Q net7 VSS VPW n18 W=720.00n L=180.00n
MM2 net5 net7 VSS VPW n18 W=0.435u L=180.00n
MM14 net_57 RDN VSS VPW n18 W=0.42u L=180.00n
MM15 net_61 net5 net_57 VPW n18 W=0.42u L=180.00n
MM17 net_45 D net_49 VPW n18 W=0.43u L=180.00n
MM18 net_49 RDN VSS VPW n18 W=0.43u L=180.00n
MM4 enn en VSS VPW n18 W=430.00n L=180.00n
MM6 en E VSS VPW n18 W=430.00n L=180.00n
.ENDS LAHRNQUHDV1
.SUBCKT LAHRNQUHDV2 D E Q RDN VDD VSS VNW VPW
MM6 en E VSS VPW n18 W=430.00n L=180.00n
MM20 net_132 en net_84 VPW n18 W=0.42u L=180.00n
MM19 net_132 enn net_80 VPW n18 W=0.43u L=180.00n
MM0 Q net_132 VSS VPW n18 W=1.44u L=180.00n
MM2 net5 net_132 VSS VPW n18 W=0.435u L=180.00n
MM18 net_76 RDN VSS VPW n18 W=0.43u L=180.00n
MM4 enn en VSS VPW n18 W=430.00n L=180.00n
MM17 net_80 D net_76 VPW n18 W=0.43u L=180.00n
MM15 net_84 net5 net_88 VPW n18 W=0.42u L=180.00n
MM14 net_88 RDN VSS VPW n18 W=0.42u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM7 en E VDD VNW p18 W=0.96u L=180.00n
MM8 net_132 RDN VDD VNW p18 W=0.73u L=180.00n
MM13 net_127 net5 VDD VNW p18 W=0.95u L=180.00n
MM11 net_132 enn net_127 VNW p18 W=0.95u L=180.00n
MM10 net_135 D VDD VNW p18 W=0.52u L=180.00n
MM9 net_132 en net_135 VNW p18 W=0.76u L=180.00n
MM3 net5 net_132 VDD VNW p18 W=0.42u L=180.00n
MM1 Q net_132 VDD VNW p18 W=2.02u L=180.00n
.ENDS LAHRNQUHDV2
.SUBCKT LAHRNQUHDV3 D E Q RDN VDD VSS VNW VPW
MM0 Q net_132 VSS VPW n18 W=2.16u L=180.00n
MM2 net5 net_132 VSS VPW n18 W=0.435u L=180.00n
MM20 net_132 en net_84 VPW n18 W=0.42u L=180.00n
MM19 net_132 enn net_80 VPW n18 W=0.43u L=180.00n
MM14 net_88 RDN VSS VPW n18 W=0.42u L=180.00n
MM15 net_84 net5 net_88 VPW n18 W=0.42u L=180.00n
MM17 net_80 D net_76 VPW n18 W=0.43u L=180.00n
MM18 net_76 RDN VSS VPW n18 W=0.49u L=180.00n
MM4 enn en VSS VPW n18 W=460.00n L=180.00n
MM6 en E VSS VPW n18 W=0.455u L=180.00n
MM1 Q net_132 VDD VNW p18 W=3.03u L=180.00n
MM3 net5 net_132 VDD VNW p18 W=0.405u L=180.00n
MM9 net_132 en net_135 VNW p18 W=0.76u L=180.00n
MM10 net_135 D VDD VNW p18 W=0.52u L=180.00n
MM11 net_132 enn net_127 VNW p18 W=0.73u L=180.00n
MM13 net_127 net5 VDD VNW p18 W=0.73u L=180.00n
MM8 net_132 RDN VDD VNW p18 W=0.73u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM7 en E VDD VNW p18 W=0.965u L=180.00n
.ENDS LAHRNQUHDV3
****Sub-Circuit for LAHSQUHDV0P7, Tue Jun 13 18:01:03 CST 2017****
.SUBCKT LAHSQUHDV0P7 D E Q SD VDD VSS VNW VPW
MM0 Q net6 VSS VPW n18 W=560.00n L=180.00n
MM2 net4 net6 VSS VPW n18 W=0.57u L=180.00n
MM4 enn en VSS VPW n18 W=460.00n L=180.00n
MM6 en E VSS VPW n18 W=0.455u L=180.00n
MM14 net_61 net4 VSS VPW n18 W=0.42u L=180.00n
MM15 net6 en net_61 VPW n18 W=0.42u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM17 net6 enn net_77 VPW n18 W=0.43u L=180.00n
MM18 net_77 D VSS VPW n18 W=0.43u L=180.00n
MM1 Q net6 VDD VNW p18 W=790.00n L=180.00n
MM3 net4 net6 VDD VNW p18 W=0.8u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM7 en E VDD VNW p18 W=0.965u L=180.00n
MM8 net_28 SD VDD VNW p18 W=0.495u L=180.00n
MM9 net_32 net4 net_28 VNW p18 W=0.495u L=180.00n
MM10 net6 enn net_32 VNW p18 W=0.495u L=180.00n
MM11 net6 en net_36 VNW p18 W=0.76u L=180.00n
MM12 net_36 D net_40 VNW p18 W=0.52u L=180.00n
MM13 net_40 SD VDD VNW p18 W=0.42u L=180.00n
.ENDS LAHSQUHDV0P7
.SUBCKT LAHSQUHDV1 D E Q SD VDD VSS VNW VPW
MM18 net_8 D VSS VPW n18 W=0.43u L=180.00n
MM17 net6 enn net_8 VPW n18 W=0.43u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM15 net6 en net_24 VPW n18 W=0.42u L=180.00n
MM14 net_24 net4 VSS VPW n18 W=0.42u L=180.00n
MM6 en E VSS VPW n18 W=0.455u L=180.00n
MM4 enn en VSS VPW n18 W=460.00n L=180.00n
MM2 net4 net6 VSS VPW n18 W=0.57u L=180.00n
MM0 Q net6 VSS VPW n18 W=720.00n L=180.00n
MM13 net_51 SD VDD VNW p18 W=0.42u L=180.00n
MM12 net_55 D net_51 VNW p18 W=0.52u L=180.00n
MM11 net6 en net_55 VNW p18 W=0.76u L=180.00n
MM10 net6 enn net_59 VNW p18 W=0.495u L=180.00n
MM9 net_59 net4 net_63 VNW p18 W=0.495u L=180.00n
MM8 net_63 SD VDD VNW p18 W=0.495u L=180.00n
MM7 en E VDD VNW p18 W=0.965u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM3 net4 net6 VDD VNW p18 W=1.01u L=180.00n
MM1 Q net6 VDD VNW p18 W=1.01u L=180.00n
.ENDS LAHSQUHDV1
.SUBCKT LAHSQUHDV2 D E Q SD VDD VSS VNW VPW
MM13 net_107 SD VDD VNW p18 W=0.425u L=180.00n
MM12 net_103 D net_107 VNW p18 W=0.52u L=180.00n
MM11 net6 en net_103 VNW p18 W=0.76u L=180.00n
MM10 net6 enn net_99 VNW p18 W=0.53u L=180.00n
MM9 net_99 net4 net_95 VNW p18 W=0.53u L=180.00n
MM8 net_95 SD VDD VNW p18 W=0.53u L=180.00n
MM7 en E VDD VNW p18 W=0.965u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM3 net4 net6 VDD VNW p18 W=1.01u L=180.00n
MM1 Q net6 VDD VNW p18 W=2.02u L=180.00n
MM18 net_144 D VSS VPW n18 W=0.43u L=180.00n
MM17 net6 enn net_144 VPW n18 W=0.43u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM15 net6 en net_128 VPW n18 W=0.42u L=180.00n
MM14 net_128 net4 VSS VPW n18 W=0.42u L=180.00n
MM6 en E VSS VPW n18 W=0.455u L=180.00n
MM4 enn en VSS VPW n18 W=460.00n L=180.00n
MM2 net4 net6 VSS VPW n18 W=0.72u L=180.00n
MM0 Q net6 VSS VPW n18 W=1.44u L=180.00n
.ENDS LAHSQUHDV2
.SUBCKT LAHSQUHDV3 D E Q SD VDD VSS VNW VPW
MM13 net_107 SD VDD VNW p18 W=0.425u L=180.00n
MM12 net_103 D net_107 VNW p18 W=0.52u L=180.00n
MM11 net6 en net_103 VNW p18 W=0.76u L=180.00n
MM10 net6 enn net_99 VNW p18 W=0.53u L=180.00n
MM9 net_99 net4 net_95 VNW p18 W=0.53u L=180.00n
MM8 net_95 SD VDD VNW p18 W=0.53u L=180.00n
MM7 en E VDD VNW p18 W=0.965u L=180.00n
MM5 enn en VDD VNW p18 W=0.89u L=180.00n
MM3 net4 net6 VDD VNW p18 W=1.01u L=180.00n
MM1 Q net6 VDD VNW p18 W=3.03u L=180.00n
MM17 net6 enn net_144 VPW n18 W=0.43u L=180.00n
MM18 net_144 D VSS VPW n18 W=0.43u L=180.00n
MM15 net6 en net_128 VPW n18 W=0.42u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM6 en E VSS VPW n18 W=0.455u L=180.00n
MM14 net_128 net4 VSS VPW n18 W=0.42u L=180.00n
MM2 net4 net6 VSS VPW n18 W=0.72u L=180.00n
MM4 enn en VSS VPW n18 W=460.00n L=180.00n
MM0 Q net6 VSS VPW n18 W=2.16u L=180.00n
.ENDS LAHSQUHDV3
.SUBCKT LALQUHDV0P7 D EN Q VDD VSS VNW VPW
MM9 cn EN VSS VPW n18 W=430.00n L=180.00n
MM6 c cn VSS VPW n18 W=670.00n L=180.00n
MM4 net24 net28 VSS VPW n18 W=0.435u L=180.00n
MM0 net32 D VSS VPW n18 W=0.42u L=180.00n
MM1 net28 cn net32 VPW n18 W=0.42u L=180.00n
MM25 Q net28 VSS VPW n18 W=0.565u L=180.00n
MM22 net16 net24 VSS VPW n18 W=0.42u L=180.00n
MM23 net28 c net16 VPW n18 W=0.42u L=180.00n
MM8 cn EN VDD VNW p18 W=0.59u L=180.00n
MM7 c cn VDD VNW p18 W=0.95u L=180.00n
MM5 net24 net28 VDD VNW p18 W=0.59u L=180.00n
MM3 net67 D VDD VNW p18 W=0.575u L=180.00n
MM2 net28 c net67 VNW p18 W=0.59u L=180.00n
MM24 Q net28 VDD VNW p18 W=0.795u L=180.00n
MM20 net28 cn net51 VNW p18 W=0.585u L=180.00n
MM21 net51 net24 VDD VNW p18 W=0.585u L=180.00n
.ENDS LALQUHDV0P7
.SUBCKT LALQUHDV1 D EN Q VDD VSS VNW VPW
MM0 net36 D VSS VPW n18 W=430.00n L=180.00n
MM1 net40 cn net36 VPW n18 W=430.00n L=180.00n
MM4 net44 net40 VSS VPW n18 W=0.44u L=180.00n
MM23 net40 c net52 VPW n18 W=430.00n L=180.00n
MM22 net52 net44 VSS VPW n18 W=430.00n L=180.00n
MM25 Q net40 VSS VPW n18 W=720.00n L=180.00n
MM6 c cn VSS VPW n18 W=0.67u L=180.00n
MM9 cn EN VSS VPW n18 W=430.00n L=180.00n
MM2 net40 c net7 VNW p18 W=0.59u L=180.00n
MM3 net7 D VDD VNW p18 W=0.59u L=180.00n
MM5 net44 net40 VDD VNW p18 W=0.585u L=180.00n
MM21 net23 net44 VDD VNW p18 W=0.59u L=180.00n
MM20 net40 cn net23 VNW p18 W=0.59u L=180.00n
MM24 Q net40 VDD VNW p18 W=1.01u L=180.00n
MM7 c cn VDD VNW p18 W=1.01u L=180.00n
MM8 cn EN VDD VNW p18 W=0.59u L=180.00n
.ENDS LALQUHDV1
.SUBCKT LALQUHDV2 D EN Q VDD VSS VNW VPW
MM0 net36 D VSS VPW n18 W=0.635u L=180.00n
MM1 net40 cn net36 VPW n18 W=0.635u L=180.00n
MM4 net44 net40 VSS VPW n18 W=0.435u L=180.00n
MM23 net40 c net52 VPW n18 W=0.435u L=180.00n
MM22 net52 net44 VSS VPW n18 W=0.435u L=180.00n
MM25 Q net40 VSS VPW n18 W=1.44u L=180.00n
MM6 c cn VSS VPW n18 W=0.67u L=180.00n
MM9 cn EN VSS VPW n18 W=430.00n L=180.00n
MM2 net40 c net7 VNW p18 W=0.945u L=180.00n
MM3 net7 D VDD VNW p18 W=0.945u L=180.00n
MM5 net44 net40 VDD VNW p18 W=0.585u L=180.00n
MM21 net23 net44 VDD VNW p18 W=0.585u L=180.00n
MM20 net40 cn net23 VNW p18 W=0.585u L=180.00n
MM24 Q net40 VDD VNW p18 W=2.02u L=180.00n
MM7 c cn VDD VNW p18 W=1.01u L=180.00n
MM8 cn EN VDD VNW p18 W=0.59u L=180.00n
.ENDS LALQUHDV2
.SUBCKT LALQUHDV3 D EN Q VDD VSS VNW VPW
MM9 cn EN VSS VPW n18 W=430.00n L=180.00n
MM6 c cn VSS VPW n18 W=0.67u L=180.00n
MM25 Q net28 VSS VPW n18 W=2.16u L=180.00n
MM22 net16 net24 VSS VPW n18 W=0.435u L=180.00n
MM23 net28 c net16 VPW n18 W=0.435u L=180.00n
MM4 net24 net28 VSS VPW n18 W=0.435u L=180.00n
MM1 net28 cn net32 VPW n18 W=0.635u L=180.00n
MM0 net32 D VSS VPW n18 W=0.635u L=180.00n
MM8 cn EN VDD VNW p18 W=0.59u L=180.00n
MM7 c cn VDD VNW p18 W=1.01u L=180.00n
MM24 Q net28 VDD VNW p18 W=3.03u L=180.00n
MM20 net28 cn net51 VNW p18 W=0.585u L=180.00n
MM21 net51 net24 VDD VNW p18 W=0.585u L=180.00n
MM5 net24 net28 VDD VNW p18 W=0.585u L=180.00n
MM3 net67 D VDD VNW p18 W=0.945u L=180.00n
MM2 net28 c net67 VNW p18 W=0.945u L=180.00n
.ENDS LALQUHDV3
.SUBCKT LALRNQUHDV0P7 D EN Q RDN VDD VSS VNW VPW
MM6 c EN VSS VPW n18 W=430.00n L=180.00n
MM4 cn c VSS VPW n18 W=430.00n L=180.00n
MM18 net_13 RDN VSS VPW n18 W=0.43u L=180.00n
MM17 net_17 D net_13 VPW n18 W=0.43u L=180.00n
MM15 net_21 net5 net_25 VPW n18 W=0.42u L=180.00n
MM14 net_25 RDN VSS VPW n18 W=0.42u L=180.00n
MM19 net_69 c net_17 VPW n18 W=0.43u L=180.00n
MM20 net_69 cn net_21 VPW n18 W=0.42u L=180.00n
MM2 net5 net_69 VSS VPW n18 W=0.435u L=180.00n
MM0 Q net_69 VSS VPW n18 W=560.00n L=180.00n
MM7 c EN VDD VNW p18 W=0.96u L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM8 net_69 RDN VDD VNW p18 W=0.505u L=180.00n
MM13 net_64 net5 VDD VNW p18 W=890.00n L=180.00n
MM11 net_69 c net_64 VNW p18 W=890.00n L=180.00n
MM10 net_72 D VDD VNW p18 W=0.52u L=180.00n
MM9 net_69 cn net_72 VNW p18 W=520.00n L=180.00n
MM3 net5 net_69 VDD VNW p18 W=490.0n L=180.00n
MM1 Q net_69 VDD VNW p18 W=0.8u L=180.00n
.ENDS LALRNQUHDV0P7
.SUBCKT LALRNQUHDV1 D EN Q RDN VDD VSS VNW VPW
MM20 net7 cn net_61 VPW n18 W=0.42u L=180.00n
MM19 net7 c net_45 VPW n18 W=0.43u L=180.00n
MM0 Q net7 VSS VPW n18 W=720.00n L=180.00n
MM2 net5 net7 VSS VPW n18 W=0.435u L=180.00n
MM14 net_57 RDN VSS VPW n18 W=0.42u L=180.00n
MM15 net_61 net5 net_57 VPW n18 W=0.42u L=180.00n
MM17 net_45 D net_49 VPW n18 W=0.43u L=180.00n
MM18 net_49 RDN VSS VPW n18 W=0.43u L=180.00n
MM4 cn c VSS VPW n18 W=430.00n L=180.00n
MM6 c EN VSS VPW n18 W=430.00n L=180.00n
MM1 Q net7 VDD VNW p18 W=1.01u L=180.00n
MM3 net5 net7 VDD VNW p18 W=490.0n L=180.00n
MM8 net7 RDN VDD VNW p18 W=0.505u L=180.00n
MM9 net7 cn net_16 VNW p18 W=520.00n L=180.00n
MM10 net_16 D VDD VNW p18 W=0.52u L=180.00n
MM11 net7 c net_20 VNW p18 W=890.00n L=180.00n
MM13 net_20 net5 VDD VNW p18 W=890.00n L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM7 c EN VDD VNW p18 W=0.96u L=180.00n
.ENDS LALRNQUHDV1
.SUBCKT LALRNQUHDV2 D EN Q RDN VDD VSS VNW VPW
MM6 c EN VSS VPW n18 W=430.00n L=180.00n
MM20 net_132 cn net_84 VPW n18 W=0.42u L=180.00n
MM19 net_132 c net_80 VPW n18 W=0.43u L=180.00n
MM0 Q net_132 VSS VPW n18 W=1.44u L=180.00n
MM2 net5 net_132 VSS VPW n18 W=0.435u L=180.00n
MM18 net_76 RDN VSS VPW n18 W=0.43u L=180.00n
MM4 cn c VSS VPW n18 W=430.00n L=180.00n
MM17 net_80 D net_76 VPW n18 W=0.43u L=180.00n
MM15 net_84 net5 net_88 VPW n18 W=0.42u L=180.00n
MM14 net_88 RDN VSS VPW n18 W=0.42u L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM7 c EN VDD VNW p18 W=0.96u L=180.00n
MM8 net_132 RDN VDD VNW p18 W=0.73u L=180.00n
MM13 net_127 net5 VDD VNW p18 W=890.00n L=180.00n
MM11 net_132 c net_127 VNW p18 W=890.00n L=180.00n
MM10 net_135 D VDD VNW p18 W=0.52u L=180.00n
MM9 net_132 cn net_135 VNW p18 W=520.00n L=180.00n
MM3 net5 net_132 VDD VNW p18 W=0.42u L=180.00n
MM1 Q net_132 VDD VNW p18 W=2.02u L=180.00n
.ENDS LALRNQUHDV2
.SUBCKT LALRNQUHDV3 D EN Q RDN VDD VSS VNW VPW
MM0 Q net_132 VSS VPW n18 W=2.16u L=180.00n
MM2 net5 net_132 VSS VPW n18 W=0.435u L=180.00n
MM20 net_132 cn net_84 VPW n18 W=0.42u L=180.00n
MM19 net_132 c net_80 VPW n18 W=0.43u L=180.00n
MM14 net_88 RDN VSS VPW n18 W=0.42u L=180.00n
MM15 net_84 net5 net_88 VPW n18 W=0.42u L=180.00n
MM17 net_80 D net_76 VPW n18 W=0.43u L=180.00n
MM18 net_76 RDN VSS VPW n18 W=0.49u L=180.00n
MM4 cn c VSS VPW n18 W=460.00n L=180.00n
MM6 c EN VSS VPW n18 W=0.455u L=180.00n
MM1 Q net_132 VDD VNW p18 W=3.03u L=180.00n
MM3 net5 net_132 VDD VNW p18 W=0.405u L=180.00n
MM9 net_132 cn net_135 VNW p18 W=520.00n L=180.00n
MM10 net_135 D VDD VNW p18 W=0.52u L=180.00n
MM11 net_132 c net_127 VNW p18 W=0.73u L=180.00n
MM13 net_127 net5 VDD VNW p18 W=0.73u L=180.00n
MM8 net_132 RDN VDD VNW p18 W=0.73u L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM7 c EN VDD VNW p18 W=0.965u L=180.00n
.ENDS LALRNQUHDV3
****Sub-Circuit for LALSQUHDV0P7, Tue Jun 13 18:01:03 CST 2017****
.SUBCKT LALSQUHDV0P7 D EN Q SD VDD VSS VNW VPW
MM0 Q net6 VSS VPW n18 W=560.00n L=180.00n
MM2 net4 net6 VSS VPW n18 W=0.57u L=180.00n
MM4 cn c VSS VPW n18 W=460.00n L=180.00n
MM6 c EN VSS VPW n18 W=0.455u L=180.00n
MM14 net_61 net4 VSS VPW n18 W=0.42u L=180.00n
MM15 net6 cn net_61 VPW n18 W=0.42u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM17 net6 c net_77 VPW n18 W=0.43u L=180.00n
MM18 net_77 D VSS VPW n18 W=0.43u L=180.00n
MM1 Q net6 VDD VNW p18 W=790.00n L=180.00n
MM3 net4 net6 VDD VNW p18 W=0.8u L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM7 c EN VDD VNW p18 W=0.965u L=180.00n
MM8 net_28 SD VDD VNW p18 W=0.495u L=180.00n
MM9 net_32 net4 net_28 VNW p18 W=435.00n L=180.00n
MM10 net6 c net_32 VNW p18 W=435.00n L=180.00n
MM11 net6 cn net_36 VNW p18 W=520.00n L=180.00n
MM12 net_36 D net_40 VNW p18 W=0.52u L=180.00n
MM13 net_40 SD VDD VNW p18 W=0.42u L=180.00n
.ENDS LALSQUHDV0P7
.SUBCKT LALSQUHDV1 D EN Q SD VDD VSS VNW VPW
MM18 net_8 D VSS VPW n18 W=0.43u L=180.00n
MM17 net6 c net_8 VPW n18 W=0.43u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM15 net6 cn net_24 VPW n18 W=0.42u L=180.00n
MM14 net_24 net4 VSS VPW n18 W=0.42u L=180.00n
MM6 c EN VSS VPW n18 W=0.455u L=180.00n
MM4 cn c VSS VPW n18 W=460.00n L=180.00n
MM2 net4 net6 VSS VPW n18 W=570.00n L=180.00n
MM0 Q net6 VSS VPW n18 W=720.00n L=180.00n
MM13 net_51 SD VDD VNW p18 W=0.42u L=180.00n
MM12 net_55 D net_51 VNW p18 W=0.52u L=180.00n
MM11 net6 cn net_55 VNW p18 W=520.00n L=180.00n
MM10 net6 c net_59 VNW p18 W=435.00n L=180.00n
MM9 net_59 net4 net_63 VNW p18 W=435.00n L=180.00n
MM8 net_63 SD VDD VNW p18 W=0.495u L=180.00n
MM7 c EN VDD VNW p18 W=0.965u L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM3 net4 net6 VDD VNW p18 W=1.01u L=180.00n
MM1 Q net6 VDD VNW p18 W=1.01u L=180.00n
.ENDS LALSQUHDV1
.SUBCKT LALSQUHDV2 D EN Q SD VDD VSS VNW VPW
MM18 net_144 D VSS VPW n18 W=0.43u L=180.00n
MM17 net6 c net_144 VPW n18 W=0.43u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM15 net6 cn net_128 VPW n18 W=0.42u L=180.00n
MM14 net_128 net4 VSS VPW n18 W=0.42u L=180.00n
MM6 c EN VSS VPW n18 W=0.455u L=180.00n
MM4 cn c VSS VPW n18 W=460.00n L=180.00n
MM2 net4 net6 VSS VPW n18 W=0.72u L=180.00n
MM0 Q net6 VSS VPW n18 W=1.44u L=180.00n
MM13 net_107 SD VDD VNW p18 W=0.425u L=180.00n
MM12 net_103 D net_107 VNW p18 W=0.52u L=180.00n
MM11 net6 cn net_103 VNW p18 W=520.00n L=180.00n
MM10 net6 c net_99 VNW p18 W=470.00n L=180.00n
MM9 net_99 net4 net_95 VNW p18 W=470.00n L=180.00n
MM8 net_95 SD VDD VNW p18 W=0.53u L=180.00n
MM7 c EN VDD VNW p18 W=0.965u L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM3 net4 net6 VDD VNW p18 W=1.01u L=180.00n
MM1 Q net6 VDD VNW p18 W=2.02u L=180.00n
.ENDS LALSQUHDV2
.SUBCKT LALSQUHDV3 D EN Q SD VDD VSS VNW VPW
MM17 net6 c net_144 VPW n18 W=0.43u L=180.00n
MM18 net_144 D VSS VPW n18 W=0.43u L=180.00n
MM15 net6 cn net_128 VPW n18 W=0.42u L=180.00n
MM16 net6 SD VSS VPW n18 W=0.57u L=180.00n
MM6 c EN VSS VPW n18 W=0.455u L=180.00n
MM14 net_128 net4 VSS VPW n18 W=0.42u L=180.00n
MM2 net4 net6 VSS VPW n18 W=0.72u L=180.00n
MM4 cn c VSS VPW n18 W=460.00n L=180.00n
MM0 Q net6 VSS VPW n18 W=2.16u L=180.00n
MM13 net_107 SD VDD VNW p18 W=0.425u L=180.00n
MM12 net_103 D net_107 VNW p18 W=0.52u L=180.00n
MM11 net6 cn net_103 VNW p18 W=520.00n L=180.00n
MM10 net6 c net_99 VNW p18 W=470.00n L=180.00n
MM9 net_99 net4 net_95 VNW p18 W=470.00n L=180.00n
MM8 net_95 SD VDD VNW p18 W=0.53u L=180.00n
MM7 c EN VDD VNW p18 W=0.965u L=180.00n
MM5 cn c VDD VNW p18 W=0.89u L=180.00n
MM3 net4 net6 VDD VNW p18 W=1.01u L=180.00n
MM1 Q net6 VDD VNW p18 W=3.03u L=180.00n
.ENDS LALSQUHDV3
****Sub-Circuit for MAJ23UHDV0P4, Thu Jun  8 09:49:35 CST 2017****
.SUBCKT MAJ23UHDV0P4 A1 A2 A3 Z VDD VSS VNW VPW
MM9 net13 A2 VSS VPW n18 W=280.00n L=180.00n
MM8 net21 A1 net13 VPW n18 W=280.00n L=180.00n
MM5 net9 A2 VSS VPW n18 W=280.00n L=180.00n
MM2 net9 A1 VSS VPW n18 W=280.00n L=180.00n
MM4 net21 A3 net9 VPW n18 W=280.00n L=180.00n
MM11 Z net21 VSS VPW n18 W=270.00n L=180.00n
MM10 Z net21 VDD VNW p18 W=490.00n L=180.00n
MM7 net21 A1 net32 VNW p18 W=490.00n L=180.00n
MM6 net32 A2 VDD VNW p18 W=490.00n L=180.00n
MM3 net21 A3 net49 VNW p18 W=490.00n L=180.00n
MM0 net49 A2 VDD VNW p18 W=490.00n L=180.00n
MM1 net49 A1 VDD VNW p18 W=490.00n L=180.00n
.ENDS MAJ23UHDV0P4
****Sub-Circuit for MAJ23UHDV0P7, Thu Jun  8 09:49:35 CST 2017****
.SUBCKT MAJ23UHDV0P7 A1 A2 A3 Z VDD VSS VNW VPW
MM9 net13 A2 VSS VPW n18 W=430.00n L=180.00n
MM8 net21 A1 net13 VPW n18 W=430.00n L=180.00n
MM5 net9 A2 VSS VPW n18 W=370.00n L=180.00n
MM2 net9 A1 VSS VPW n18 W=430.00n L=180.00n
MM4 net21 A3 net9 VPW n18 W=370.00n L=180.00n
MM11 Z net21 VSS VPW n18 W=560.00n L=180.00n
MM10 Z net21 VDD VNW p18 W=790.0n L=180.00n
MM7 net21 A1 net32 VNW p18 W=500.00n L=180.00n
MM6 net32 A2 VDD VNW p18 W=500.00n L=180.00n
MM3 net21 A3 net49 VNW p18 W=500.00n L=180.00n
MM0 net49 A2 VDD VNW p18 W=500.00n L=180.00n
MM1 net49 A1 VDD VNW p18 W=500.00n L=180.00n
.ENDS MAJ23UHDV0P7
****Sub-Circuit for MAJ23UHDV1, Thu Jun  8 09:49:35 CST 2017****
.SUBCKT MAJ23UHDV1 A1 A2 A3 Z VDD VSS VNW VPW
MM9 net13 A2 VSS VPW n18 W=430.00n L=180.00n
MM8 net21 A1 net13 VPW n18 W=430.00n L=180.00n
MM5 net9 A2 VSS VPW n18 W=370.00n L=180.00n
MM2 net9 A1 VSS VPW n18 W=430.00n L=180.00n
MM4 net21 A3 net9 VPW n18 W=370.00n L=180.00n
MM11 Z net21 VSS VPW n18 W=720.00n L=180.00n
MM10 Z net21 VDD VNW p18 W=1.01u L=180.00n
MM7 net21 A1 net32 VNW p18 W=580.00n L=180.00n
MM6 net32 A2 VDD VNW p18 W=580.00n L=180.00n
MM3 net21 A3 net49 VNW p18 W=510.00n L=180.00n
MM0 net49 A2 VDD VNW p18 W=510.00n L=180.00n
MM1 net49 A1 VDD VNW p18 W=580.00n L=180.00n
.ENDS MAJ23UHDV1
****Sub-Circuit for MAJ23UHDV2, Thu Jun  8 09:49:35 CST 2017****
.SUBCKT MAJ23UHDV2 A1 A2 A3 Z VDD VSS VNW VPW
MM9 net13 A2 VSS VPW n18 W=630.00n L=180.00n
MM8 net21 A1 net13 VPW n18 W=630.00n L=180.00n
MM5 net9 A2 VSS VPW n18 W=630.00n L=180.00n
MM2 net9 A1 VSS VPW n18 W=630.00n L=180.00n
MM4 net21 A3 net9 VPW n18 W=630.00n L=180.00n
MM11 Z net21 VSS VPW n18 W=1.44u L=180.00n
MM10 Z net21 VDD VNW p18 W=2.02u L=180.00n
MM7 net21 A1 net32 VNW p18 W=950.00n L=180.00n
MM6 net32 A2 VDD VNW p18 W=950.00n L=180.00n
MM3 net21 A3 net49 VNW p18 W=950.00n L=180.00n
MM0 net49 A2 VDD VNW p18 W=855.00n L=180.00n
MM1 net49 A1 VDD VNW p18 W=950.00n L=180.00n
.ENDS MAJ23UHDV2
****Sub-Circuit for MAJ23UHDV3, Thu Jun  8 09:49:35 CST 2017****
.SUBCKT MAJ23UHDV3 A1 A2 A3 Z VDD VSS VNW VPW
MM9 net13 A2 VSS VPW n18 W=720.00n L=180.00n
MM8 net21 A1 net13 VPW n18 W=720.00n L=180.00n
MM5 net9 A2 VSS VPW n18 W=720.00n L=180.00n
MM2 net9 A1 VSS VPW n18 W=720.00n L=180.00n
MM4 net21 A3 net9 VPW n18 W=720.00n L=180.00n
MM11 Z net21 VSS VPW n18 W=2.16u L=180.00n
MM10 Z net21 VDD VNW p18 W=3.03u L=180.00n
MM7 net21 A1 net32 VNW p18 W=1.01u L=180.00n
MM6 net32 A2 VDD VNW p18 W=1.01u L=180.00n
MM3 net21 A3 net49 VNW p18 W=1.01u L=180.00n
MM0 net49 A2 VDD VNW p18 W=915.00n L=180.00n
MM1 net49 A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS MAJ23UHDV3
****Sub-Circuit for MAOI222UHDV0P4, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MAOI222UHDV0P4 A B C ZN VDD VSS VNW VPW
MMN1 net6 B VSS VPW n18 W=280.00n L=180.00n
MM4 ZN A net5 VPW n18 W=280.00n L=180.00n
MM1 ZN A net6 VPW n18 W=280.00n L=180.00n
MM9 net5 C VSS VPW n18 W=280.00n L=180.00n
MM10 net4 C VSS VPW n18 W=280.00n L=180.00n
MM6 ZN B net4 VPW n18 W=280.00n L=180.00n
MMP1 ZN A net2 VNW p18 W=490.00n L=180.00n
MM0 net2 A net1 VNW p18 W=490.00n L=180.00n
MM5 net1 C VDD VNW p18 W=490.00n L=180.00n
MM7 net1 B VDD VNW p18 W=490.00n L=180.00n
MM11 ZN B net2 VNW p18 W=490.00n L=180.00n
MM8 net2 C net1 VNW p18 W=490.00n L=180.00n
.ENDS MAOI222UHDV0P4
****Sub-Circuit for MAOI222UHDV0P7, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MAOI222UHDV0P7 A B C ZN VDD VSS VNW VPW
MMN1 net6 B VSS VPW n18 W=560.00n L=180.00n
MM4 ZN A net5 VPW n18 W=560.00n L=180.00n
MM1 ZN A net6 VPW n18 W=560.00n L=180.00n
MM9 net5 C VSS VPW n18 W=560.00n L=180.00n
MM10 net4 C VSS VPW n18 W=560.00n L=180.00n
MM6 ZN B net4 VPW n18 W=560.00n L=180.00n
MMP1 ZN A net2 VNW p18 W=790.00n L=180.00n
MM0 net2 A net1 VNW p18 W=790.00n L=180.00n
MM5 net1 C VDD VNW p18 W=790.00n L=180.00n
MM7 net1 B VDD VNW p18 W=790.00n L=180.00n
MM11 ZN B net2 VNW p18 W=790.00n L=180.00n
MM8 net2 C net1 VNW p18 W=790.00n L=180.00n
.ENDS MAOI222UHDV0P7
****Sub-Circuit for MAOI222UHDV1, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MAOI222UHDV1 A B C ZN VDD VSS VNW VPW
MMN1 net6 B VSS VPW n18 W=720.00n L=180.00n
MM4 ZN A net5 VPW n18 W=720.00n L=180.00n
MM1 ZN A net6 VPW n18 W=720.00n L=180.00n
MM9 net5 C VSS VPW n18 W=720.00n L=180.00n
MM10 net4 C VSS VPW n18 W=720.00n L=180.00n
MM6 ZN B net4 VPW n18 W=720.00n L=180.00n
MMP1 ZN A net2 VNW p18 W=975.00n L=180.00n
MM0 net2 A net1 VNW p18 W=975.00n L=180.00n
MM5 net1 C VDD VNW p18 W=1.01u L=180.00n
MM7 net1 B VDD VNW p18 W=1.01u L=180.00n
MM11 ZN B net2 VNW p18 W=1.01u L=180.00n
MM8 net2 C net1 VNW p18 W=975.00n L=180.00n
.ENDS MAOI222UHDV1
****Sub-Circuit for MAOI222UHDV2, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MAOI222UHDV2 A B C ZN VDD VSS VNW VPW
MMN1 net6 B VSS VPW n18 W=1.44u L=180.00n
MM4 ZN A net5 VPW n18 W=620.00n L=180.00n
MM1 ZN A net6 VPW n18 W=1.44u L=180.00n
MM9 net5 C VSS VPW n18 W=1.42u L=180.00n
MM10 net4 C VSS VPW n18 W=1.44u L=180.00n
MM6 ZN B net4 VPW n18 W=1.44u L=180.00n
MMP1 ZN A net2 VNW p18 W=1.985u L=180.00n
MM0 net2 A net1 VNW p18 W=2.02u L=180.00n
MM5 net1 C VDD VNW p18 W=2.02u L=180.00n
MM7 net1 B VDD VNW p18 W=1.95u L=180.00n
MM11 ZN B net2 VNW p18 W=1.985u L=180.00n
MM8 net2 C net1 VNW p18 W=2.02u L=180.00n
.ENDS MAOI222UHDV2
****Sub-Circuit for MAOI222UHDV3, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MAOI222UHDV3 A B C ZN VDD VSS VNW VPW
MMN1 net6 B VSS VPW n18 W=2.16u L=180.00n
MM4 ZN A net5 VPW n18 W=1.3u L=180.00n
MM1 ZN A net6 VPW n18 W=2.16u L=180.00n
MM9 net5 C VSS VPW n18 W=2.04u L=180.00n
MM10 net4 C VSS VPW n18 W=2.16u L=180.00n
MM6 ZN B net4 VPW n18 W=2.16u L=180.00n
MMP1 ZN A net2 VNW p18 W=2.925u L=180.00n
MM0 net2 A net1 VNW p18 W=2.925u L=180.00n
MM5 net1 C VDD VNW p18 W=2.96u L=180.00n
MM7 net1 B VDD VNW p18 W=3.03u L=180.00n
MM11 ZN B net2 VNW p18 W=3.03u L=180.00n
MM8 net2 C net1 VNW p18 W=2.96u L=180.00n
.ENDS MAOI222UHDV3
****Sub-Circuit for MOAI222UHDV0P4, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MOAI222UHDV0P4 A B C ZN VDD VSS VNW VPW
MM5 ZN B net_48 VPW n18 W=280.00n L=180.00n
MM4 ZN A net_48 VPW n18 W=280.00n L=180.00n
MM1 net_40 C VSS VPW n18 W=280.00n L=180.00n
MM0 net_40 B VSS VPW n18 W=280.00n L=180.00n
MM3 net_48 C net_40 VPW n18 W=280.00n L=180.00n
MM2 net_48 A net_40 VPW n18 W=280.00n L=180.00n
MM10 net_87 C VDD VNW p18 W=490.00n L=180.00n
MM7 ZN A net_87 VNW p18 W=490.00n L=180.00n
MM11 net_91 C VDD VNW p18 W=490.00n L=180.00n
MM8 ZN B net_91 VNW p18 W=490.00n L=180.00n
MM6 ZN A net_99 VNW p18 W=490.00n L=180.00n
MM9 net_99 B VDD VNW p18 W=490.00n L=180.00n
.ENDS MOAI222UHDV0P4
****Sub-Circuit for MOAI222UHDV0P7, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MOAI222UHDV0P7 A B C ZN VDD VSS VNW VPW
MM5 ZN B net_48 VPW n18 W=560.00n L=180.00n
MM4 ZN A net_48 VPW n18 W=560.00n L=180.00n
MM1 net_40 C VSS VPW n18 W=560.00n L=180.00n
MM0 net_40 B VSS VPW n18 W=560.00n L=180.00n
MM3 net_48 C net_40 VPW n18 W=560.00n L=180.00n
MM2 net_48 A net_40 VPW n18 W=560.00n L=180.00n
MM10 net_87 C VDD VNW p18 W=770.00n L=180.00n
MM7 ZN A net_87 VNW p18 W=770.00n L=180.00n
MM11 net_91 C VDD VNW p18 W=790.00n L=180.00n
MM8 ZN B net_91 VNW p18 W=790.00n L=180.00n
MM6 ZN A net_99 VNW p18 W=770.00n L=180.00n
MM9 net_99 B VDD VNW p18 W=770.00n L=180.00n
.ENDS MOAI222UHDV0P7
****Sub-Circuit for MOAI222UHDV1, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MOAI222UHDV1 A B C ZN VDD VSS VNW VPW
MM5 ZN B net_48 VPW n18 W=720.00n L=180.00n
MM4 ZN A net_48 VPW n18 W=720.00n L=180.00n
MM1 net_40 C VSS VPW n18 W=720.00n L=180.00n
MM0 net_40 B VSS VPW n18 W=720.00n L=180.00n
MM3 net_48 C net_40 VPW n18 W=720.00n L=180.00n
MM2 net_48 A net_40 VPW n18 W=720.00n L=180.00n
MM10 net_87 C VDD VNW p18 W=770.00n L=180.00n
MM7 ZN A net_87 VNW p18 W=770.00n L=180.00n
MM11 net_91 C VDD VNW p18 W=1.01u L=180.00n
MM8 ZN B net_91 VNW p18 W=1.01u L=180.00n
MM6 ZN A net_99 VNW p18 W=770.00n L=180.00n
MM9 net_99 B VDD VNW p18 W=770.00n L=180.00n
.ENDS MOAI222UHDV1
****Sub-Circuit for MOAI222UHDV2, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MOAI222UHDV2 A B C ZN VDD VSS VNW VPW
MM5 ZN B net_48 VPW n18 W=1.44u L=180.00n
MM4 ZN A net_48 VPW n18 W=1.44u L=180.00n
MM1 net_40 C VSS VPW n18 W=1.44u L=180.00n
MM0 net_40 B VSS VPW n18 W=1.44u L=180.00n
MM3 net_48 C net_40 VPW n18 W=1.44u L=180.00n
MM2 net_48 A net_40 VPW n18 W=1.44u L=180.00n
MM10 net_87 C VDD VNW p18 W=2.005u L=180.00n
MM7 ZN A net_87 VNW p18 W=1.62u L=180.00n
MM11 net_91 C VDD VNW p18 W=1.78u L=180.00n
MM8 ZN B net_91 VNW p18 W=1.78u L=180.00n
MM6 ZN A net_99 VNW p18 W=1.54u L=180.00n
MM9 net_99 B VDD VNW p18 W=1.54u L=180.00n
.ENDS MOAI222UHDV2
****Sub-Circuit for MOAI222UHDV3, Tue Jun  6 17:50:08 CST 2017****
.SUBCKT MOAI222UHDV3 A B C ZN VDD VSS VNW VPW
MM5 ZN B net_48 VPW n18 W=2.16u L=180.00n
MM4 ZN A net_48 VPW n18 W=2.16u L=180.00n
MM1 net_40 C VSS VPW n18 W=2.16u L=180.00n
MM0 net_40 B VSS VPW n18 W=2.16u L=180.00n
MM3 net_48 C net_40 VPW n18 W=2.16u L=180.00n
MM2 net_48 A net_40 VPW n18 W=2.16u L=180.00n
MM10 net_87 C VDD VNW p18 W=2.65u L=180.00n
MM7 ZN A net_87 VNW p18 W=2.47u L=180.00n
MM11 net_91 C VDD VNW p18 W=2.55u L=180.00n
MM8 ZN B net_91 VNW p18 W=3.03u L=180.00n
MM6 ZN A net_99 VNW p18 W=2.31u L=180.00n
MM9 net_99 B VDD VNW p18 W=2.61u L=180.00n
.ENDS MOAI222UHDV3
.SUBCKT MUX2NUHDV0P4 I0 I1 S ZN VDD VSS VNW VPW
MM10 SN S VDD VNW p18 W=490.0n L=180.00n
MM1 ZN S net12 VNW p18 W=490.0n L=180.00n
MM2 net12 I0 VDD VNW p18 W=490.0n L=180.00n
MM6 net24 I1 VDD VNW p18 W=490.0n L=180.00n
MM7 ZN SN net24 VNW p18 W=490.0n L=180.00n
MM11 SN S VSS VPW n18 W=0.28u L=180.00n
MM0 ZN SN net33 VPW n18 W=0.28u L=180.00n
MM3 net33 I0 VSS VPW n18 W=0.28u L=180.00n
MM4 net37 I1 VSS VPW n18 W=0.28u L=180.00n
MM5 ZN S net37 VPW n18 W=0.28u L=180.00n
.ENDS MUX2NUHDV0P4
.SUBCKT MUX2NUHDV0P7 I0 I1 S ZN VDD VSS VNW VPW
MM5 ZN S net9 VPW n18 W=560.00n L=180.00n
MM4 net9 I1 VSS VPW n18 W=560.00n L=180.00n
MM3 net13 I0 VSS VPW n18 W=560.00n L=180.00n
MM0 ZN SN net13 VPW n18 W=560.00n L=180.00n
MM11 SN S VSS VPW n18 W=560.00n L=180.00n
MM7 ZN SN net28 VNW p18 W=790.0n L=180.00n
MM6 net28 I1 VDD VNW p18 W=790.0n L=180.00n
MM2 net40 I0 VDD VNW p18 W=580.00n L=180.00n
MM1 ZN S net40 VNW p18 W=790.0n L=180.00n
MM10 SN S VDD VNW p18 W=790.00n L=180.00n
.ENDS MUX2NUHDV0P7
.SUBCKT MUX2NUHDV1 I0 I1 S ZN VDD VSS VNW VPW
MM5 ZN S net9 VPW n18 W=0.42u L=180.00n
MM4 net9 I1 VSS VPW n18 W=0.37u L=180.00n
MM3 net13 I0 VSS VPW n18 W=690.00n L=180.00n
MM0 ZN SN net13 VPW n18 W=690.00n L=180.00n
MM11 SN S VSS VPW n18 W=0.66u L=180.00n
MM7 ZN SN net28 VNW p18 W=0.58u L=180.00n
MM6 net28 I1 VDD VNW p18 W=0.58u L=180.00n
MM2 net40 I0 VDD VNW p18 W=0.95u L=180.00n
MM1 ZN S net40 VNW p18 W=0.95u L=180.00n
MM10 SN S VDD VNW p18 W=0.95u L=180.00n
.ENDS MUX2NUHDV1
.SUBCKT MUX2NUHDV2 I0 I1 S ZN VDD VSS VNW VPW
MM5 ZN S net9 VPW n18 W=0.86u L=180.00n
MM4 net9 I1 VSS VPW n18 W=1.32u L=180.00n
MM3 net13 I0 VSS VPW n18 W=1.335u L=180.00n
MM0 ZN SN net13 VPW n18 W=0.615u L=180.00n
MM11 SN S VSS VPW n18 W=0.66u L=180.00n
MM7 ZN SN net28 VNW p18 W=0.95u L=180.00n
MM6 net28 I1 VDD VNW p18 W=2.02u L=180.00n
MM2 net40 I0 VDD VNW p18 W=1.9u L=180.00n
MM1 ZN S net40 VNW p18 W=0.95u L=180.00n
MM10 SN S VDD VNW p18 W=1.405u L=180.00n
.ENDS MUX2NUHDV2
.SUBCKT MUX2UHDV0P4 I0 I1 S Z VDD VSS VNW VPW
MM8 Z net35 VSS VPW n18 W=0.28u L=180.00n
MM5 net35 S net27 VPW n18 W=0.28u L=180.00n
MM4 net27 I1 VSS VPW n18 W=0.28u L=180.00n
MM3 net31 I0 VSS VPW n18 W=0.28u L=180.00n
MM0 net35 SN net31 VPW n18 W=0.28u L=180.00n
MM12 SN S VSS VPW n18 W=0.28u L=180.00n
MM9 Z net35 VDD VNW p18 W=490.0n L=180.00n
MM7 net35 SN net50 VNW p18 W=490.0n L=180.00n
MM6 net50 I1 VDD VNW p18 W=490.0n L=180.00n
MM2 net62 I0 VDD VNW p18 W=490.0n L=180.00n
MM1 net35 S net62 VNW p18 W=490.0n L=180.00n
MM13 SN S VDD VNW p18 W=490.0n L=180.00n
.ENDS MUX2UHDV0P4
.SUBCKT MUX2UHDV0P7 I0 I1 S Z VDD VSS VNW VPW
MM13 SN S VDD VNW p18 W=490.0n L=180.00n
MM1 net33 S net12 VNW p18 W=500.0n L=180.00n
MM2 net12 I0 VDD VNW p18 W=500.0n L=180.00n
MM6 net24 I1 VDD VNW p18 W=500.0n L=180.00n
MM7 net33 SN net24 VNW p18 W=500.0n L=180.00n
MM9 Z net33 VDD VNW p18 W=790.0n L=180.00n
MM12 SN S VSS VPW n18 W=430.00n L=180.00n
MM0 net33 SN net37 VPW n18 W=300.00n L=180.00n
MM3 net37 I0 VSS VPW n18 W=300.00n L=180.00n
MM4 net41 I1 VSS VPW n18 W=430.00n L=180.00n
MM5 net33 S net41 VPW n18 W=430.00n L=180.00n
MM8 Z net33 VSS VPW n18 W=560.00n L=180.00n
.ENDS MUX2UHDV0P7
.SUBCKT MUX2UHDV1 I0 I1 S Z VDD VSS VNW VPW
MM13 SN S VDD VNW p18 W=490.0n L=180.00n
MM1 net33 S net12 VNW p18 W=500.0n L=180.00n
MM2 net12 I0 VDD VNW p18 W=500.0n L=180.00n
MM6 net24 I1 VDD VNW p18 W=0.535u L=180.00n
MM7 net33 SN net24 VNW p18 W=0.535u L=180.00n
MM9 Z net33 VDD VNW p18 W=1.01u L=180.00n
MM12 SN S VSS VPW n18 W=430.00n L=180.00n
MM0 net33 SN net37 VPW n18 W=300.00n L=180.00n
MM3 net37 I0 VSS VPW n18 W=300.00n L=180.00n
MM4 net41 I1 VSS VPW n18 W=430.00n L=180.00n
MM5 net33 S net41 VPW n18 W=430.00n L=180.00n
MM8 Z net33 VSS VPW n18 W=720.00n L=180.00n
.ENDS MUX2UHDV1
.SUBCKT MUX2UHDV2 I0 I1 S Z VDD VSS VNW VPW
MM13 SN S VDD VNW p18 W=0.66u L=180.00n
MM1 net33 S net12 VNW p18 W=0.83u L=180.00n
MM2 net12 I0 VDD VNW p18 W=0.83u L=180.00n
MM6 net24 I1 VDD VNW p18 W=0.96u L=180.00n
MM7 net33 SN net24 VNW p18 W=0.96u L=180.00n
MM9 Z net33 VDD VNW p18 W=2.02u L=180.00n
MM12 SN S VSS VPW n18 W=460.00n L=180.00n
MM0 net33 SN net37 VPW n18 W=0.7u L=180.00n
MM3 net37 I0 VSS VPW n18 W=0.7u L=180.00n
MM4 net41 I1 VSS VPW n18 W=0.7u L=180.00n
MM5 net33 S net41 VPW n18 W=0.7u L=180.00n
MM8 Z net33 VSS VPW n18 W=1.44u L=180.00n
.ENDS MUX2UHDV2
.SUBCKT MUX2UHDV3 I0 I1 S Z VDD VSS VNW VPW
MM13 SN S VDD VNW p18 W=0.88u L=180.00n
MM1 net33 S net12 VNW p18 W=0.95u L=180.00n
MM2 net12 I0 VDD VNW p18 W=0.58u L=180.00n
MM6 net24 I1 VDD VNW p18 W=0.99u L=180.00n
MM7 net33 SN net24 VNW p18 W=0.99u L=180.00n
MM9 Z net33 VDD VNW p18 W=2.97u L=180.00n
MM12 SN S VSS VPW n18 W=700.00n L=180.00n
MM0 net33 SN net37 VPW n18 W=720.00n L=180.00n
MM3 net37 I0 VSS VPW n18 W=720.00n L=180.00n
MM4 net41 I1 VSS VPW n18 W=720.00n L=180.00n
MM5 net33 S net41 VPW n18 W=720.00n L=180.00n
MM8 Z net33 VSS VPW n18 W=2.16u L=180.00n
.ENDS MUX2UHDV3
.SUBCKT MUX2UHDV6 I0 I1 S Z VDD VSS VNW VPW
MM1 net29 S net8 VNW p18 W=1.9u L=180.00n
MM2 net8 I0 VDD VNW p18 W=2.02u L=180.00n
MM6 net20 I1 VDD VNW p18 W=2.02u L=180.00n
MM7 net29 SN net20 VNW p18 W=1.9u L=180.00n
MM9 Z net29 VDD VNW p18 W=6.06u L=180.00n
MM13 SN S VDD VNW p18 W=1.45u L=180.00n
MM0 net29 SN net33 VPW n18 W=1.44u L=180.00n
MM3 net33 I0 VSS VPW n18 W=1.44u L=180.00n
MM4 net37 I1 VSS VPW n18 W=1420.00n L=180.00n
MM5 net29 S net37 VPW n18 W=1.44u L=180.00n
MM8 Z net29 VSS VPW n18 W=4.32u L=180.00n
MM12 SN S VSS VPW n18 W=1050.00n L=180.00n
.ENDS MUX2UHDV6
.SUBCKT MUX3UHDV0P7 I0 I1 I2 S0 S1 Z VDD VSS VNW VPW
MM16 net086 I2 VDD VNW p18 W=0.51u L=180.00n
MM17 net0134 S1N net086 VNW p18 W=0.51u L=180.00n
MM10 S0N S0 VDD VNW p18 W=0.59u L=180.00n
MM14 net29 S1 net0134 VNW p18 W=0.51u L=180.00n
MM1 net29 S0 net8 VNW p18 W=0.51u L=180.00n
MM2 net8 I0 VDD VNW p18 W=0.51u L=180.00n
MM6 net20 I1 VDD VNW p18 W=0.51u L=180.00n
MM7 net29 S0N net20 VNW p18 W=0.51u L=180.00n
MM9 Z net0134 VDD VNW p18 W=0.8u L=180.00n
MM13 S1N S1 VDD VNW p18 W=0.5u L=180.00n
MM11 S0N S0 VSS VPW n18 W=430.00n L=180.00n
MM18 net0127 I2 VSS VPW n18 W=0.44u L=180.00n
MM19 net0134 S1 net0127 VPW n18 W=0.44u L=180.00n
MM15 net29 S1N net0134 VPW n18 W=0.44u L=180.00n
MM0 net29 S0N net33 VPW n18 W=0.44u L=180.00n
MM3 net33 I0 VSS VPW n18 W=0.44u L=180.00n
MM4 net37 I1 VSS VPW n18 W=0.35u L=180.00n
MM5 net29 S0 net37 VPW n18 W=0.35u L=180.00n
MM8 Z net0134 VSS VPW n18 W=0.57u L=180.00n
MM12 S1N S1 VSS VPW n18 W=0.44u L=180.00n
.ENDS MUX3UHDV0P7
.SUBCKT MUX3UHDV1 I0 I1 I2 S0 S1 Z VDD VSS VNW VPW
MM11 S0N S0 VSS VPW n18 W=430.00n L=180.00n
MM18 net162 I2 VSS VPW n18 W=0.44u L=180.00n
MM19 net157 S1 net162 VPW n18 W=0.44u L=180.00n
MM15 net150 S1N net157 VPW n18 W=0.44u L=180.00n
MM0 net150 S0N net146 VPW n18 W=0.44u L=180.00n
MM3 net146 I0 VSS VPW n18 W=0.44u L=180.00n
MM4 net142 I1 VSS VPW n18 W=0.35u L=180.00n
MM5 net150 S0 net142 VPW n18 W=0.35u L=180.00n
MM8 Z net157 VSS VPW n18 W=720.00n L=180.00n
MM12 S1N S1 VSS VPW n18 W=0.44u L=180.00n
MM17 net157 S1N net205 VNW p18 W=0.51u L=180.00n
MM16 net205 I2 VDD VNW p18 W=0.595u L=180.00n
MM14 net150 S1 net157 VNW p18 W=0.51u L=180.00n
MM10 S0N S0 VDD VNW p18 W=0.59u L=180.00n
MM2 net193 I0 VDD VNW p18 W=0.505u L=180.00n
MM1 net150 S0 net193 VNW p18 W=0.505u L=180.00n
MM7 net150 S0N net181 VNW p18 W=0.51u L=180.00n
MM6 net181 I1 VDD VNW p18 W=0.51u L=180.00n
MM13 S1N S1 VDD VNW p18 W=0.6u L=180.00n
MM9 Z net157 VDD VNW p18 W=1.01u L=180.00n
.ENDS MUX3UHDV1
.SUBCKT MUX3UHDV2 I0 I1 I2 S0 S1 Z VDD VSS VNW VPW
MM12 S1N S1 VSS VPW n18 W=0.44u L=180.00n
MM8 Z net34 VSS VPW n18 W=1.44u L=180.00n
MM5 net27 S0 net19 VPW n18 W=0.35u L=180.00n
MM4 net19 I1 VSS VPW n18 W=0.35u L=180.00n
MM3 net23 I0 VSS VPW n18 W=0.44u L=180.00n
MM0 net27 S0N net23 VPW n18 W=0.44u L=180.00n
MM15 net27 S1N net34 VPW n18 W=0.44u L=180.00n
MM19 net34 S1 net39 VPW n18 W=0.44u L=180.00n
MM18 net39 I2 VSS VPW n18 W=0.44u L=180.00n
MM11 S0N S0 VSS VPW n18 W=430.00n L=180.00n
MM13 S1N S1 VDD VNW p18 W=0.59u L=180.00n
MM9 Z net34 VDD VNW p18 W=2.02u L=180.00n
MM7 net27 S0N net58 VNW p18 W=0.51u L=180.00n
MM6 net58 I1 VDD VNW p18 W=0.51u L=180.00n
MM2 net70 I0 VDD VNW p18 W=0.51u L=180.00n
MM1 net27 S0 net70 VNW p18 W=0.51u L=180.00n
MM14 net27 S1 net34 VNW p18 W=0.51u L=180.00n
MM10 S0N S0 VDD VNW p18 W=0.59u L=180.00n
MM17 net34 S1N net82 VNW p18 W=0.8u L=180.00n
MM16 net82 I2 VDD VNW p18 W=0.8u L=180.00n
.ENDS MUX3UHDV2
.SUBCKT MUXINOR2UHDV0P7 EN I0 I1 S Z VDD VSS VNW VPW
MM9 Z EN VSS VPW n18 W=560.00n L=180.00n
MM8 Z net26 VSS VPW n18 W=560.00n L=180.00n
MM5 net26 S net18 VPW n18 W=430.00n L=180.00n
MM4 net18 I1 VSS VPW n18 W=430.00n L=180.00n
MM3 net22 I0 VSS VPW n18 W=430.00n L=180.00n
MM0 net26 SN net22 VPW n18 W=430.00n L=180.00n
MM11 SN S VSS VPW n18 W=430.00n L=180.00n
MM13 net41 EN VDD VNW p18 W=790.0n L=180.00n
MM12 Z net26 net41 VNW p18 W=790.0n L=180.00n
MM7 net26 SN net45 VNW p18 W=500.0n L=180.00n
MM6 net45 I1 VDD VNW p18 W=500.0n L=180.00n
MM2 net57 I0 VDD VNW p18 W=500.0n L=180.00n
MM1 net26 S net57 VNW p18 W=500.0n L=180.00n
MM10 SN S VDD VNW p18 W=490.0n L=180.00n
.ENDS MUXINOR2UHDV0P7
.SUBCKT MUXINOR2UHDV1 EN I0 I1 S Z VDD VSS VNW VPW
MM10 SN S VDD VNW p18 W=490.0n L=180.00n
MM1 net38 S net13 VNW p18 W=570.0n L=180.00n
MM2 net13 I0 VDD VNW p18 W=580.0n L=180.00n
MM6 net25 I1 VDD VNW p18 W=580.0n L=180.00n
MM7 net38 SN net25 VNW p18 W=580.0n L=180.00n
MM12 Z net38 net29 VNW p18 W=1.01u L=180.00n
MM13 net29 EN VDD VNW p18 W=1.01u L=180.00n
MM11 SN S VSS VPW n18 W=430.00n L=180.00n
MM0 net38 SN net42 VPW n18 W=430.00n L=180.00n
MM3 net42 I0 VSS VPW n18 W=430.00n L=180.00n
MM4 net46 I1 VSS VPW n18 W=430.00n L=180.00n
MM5 net38 S net46 VPW n18 W=430.00n L=180.00n
MM8 Z net38 VSS VPW n18 W=720.00n L=180.00n
MM9 Z EN VSS VPW n18 W=720.00n L=180.00n
.ENDS MUXINOR2UHDV1
.SUBCKT MUXINOR2UHDV2 EN I0 I1 S Z VDD VSS VNW VPW
MM9 Z EN VSS VPW n18 W=1.44u L=180.00n
MM8 Z net26 VSS VPW n18 W=1.44u L=180.00n
MM5 net26 S net18 VPW n18 W=430.00n L=180.00n
MM4 net18 I1 VSS VPW n18 W=430.00n L=180.00n
MM3 net22 I0 VSS VPW n18 W=430.00n L=180.00n
MM0 net26 SN net22 VPW n18 W=430.00n L=180.00n
MM11 SN S VSS VPW n18 W=430.00n L=180.00n
MM13 net41 EN VDD VNW p18 W=2.02u L=180.00n
MM12 Z net26 net41 VNW p18 W=2.02u L=180.00n
MM7 net26 SN net45 VNW p18 W=580.0n L=180.00n
MM6 net45 I1 VDD VNW p18 W=580.0n L=180.00n
MM2 net57 I0 VDD VNW p18 W=580.0n L=180.00n
MM1 net26 S net57 VNW p18 W=570.0n L=180.00n
MM10 SN S VDD VNW p18 W=490.0n L=180.00n
.ENDS MUXINOR2UHDV2
.SUBCKT NAND2UHDV0P4 A1 A2 ZN VDD VSS VNW VPW
MM2 ZN A1 VDD VNW p18 W=0.5u L=180.00n
MM0 ZN A2 VDD VNW p18 W=0.5u L=180.00n
MM1 ZN A1 net16 VPW n18 W=0.28u L=180.00n
MM3 net16 A2 VSS VPW n18 W=0.28u L=180.00n
.ENDS NAND2UHDV0P4
.SUBCKT NAND2UHDV0P7 A1 A2 ZN VDD VSS VNW VPW
MM3 net4 A2 VSS VPW n18 W=0.605u L=180.00n
MM1 ZN A1 net4 VPW n18 W=0.605u L=180.00n
MM0 ZN A2 VDD VNW p18 W=0.805u L=180.00n
MM2 ZN A1 VDD VNW p18 W=0.805u L=180.00n
.ENDS NAND2UHDV0P7
.SUBCKT NAND2UHDV1 A1 A2 ZN VDD VSS VNW VPW
MM3 net4 A2 VSS VPW n18 W=720.00n L=180.00n
MM1 ZN A1 net4 VPW n18 W=720.00n L=180.00n
MM0 ZN A2 VDD VNW p18 W=1.01u L=180.00n
MM2 ZN A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS NAND2UHDV1
.SUBCKT NAND2UHDV2 A1 A2 ZN VDD VSS VNW VPW
MM3 net4 A2 VSS VPW n18 W=1.44u L=180.00n
MM1 ZN A1 net4 VPW n18 W=1.44u L=180.00n
MM0 ZN A2 VDD VNW p18 W=2.02u L=180.00n
MM2 ZN A1 VDD VNW p18 W=2.02u L=180.00n
.ENDS NAND2UHDV2
.SUBCKT NAND2UHDV3 A1 A2 ZN VDD VSS VNW VPW
MM3 net4 A2 VSS VPW n18 W=2.16u L=180.00n
MM1 ZN A1 net4 VPW n18 W=2.16u L=180.00n
MM0 ZN A2 VDD VNW p18 W=2.995u L=180.00n
MM2 ZN A1 VDD VNW p18 W=3.03u L=180.00n
.ENDS NAND2UHDV3
.SUBCKT NAND2UHDV4 A1 A2 ZN VDD VSS VNW VPW
MM3 net4 A2 VSS VPW n18 W=2.88u L=180.00n
MM1 ZN A1 net4 VPW n18 W=2.88u L=180.00n
MM0 ZN A2 VDD VNW p18 W=4.005u L=180.00n
MM2 ZN A1 VDD VNW p18 W=4.04u L=180.00n
.ENDS NAND2UHDV4
.SUBCKT NAND2UHDV6 A1 A2 ZN VDD VSS VNW VPW
MM3 net4 A2 VSS VPW n18 W=4.32u L=180.00n
MM1 ZN A1 net4 VPW n18 W=4.32u L=180.00n
MM0 ZN A2 VDD VNW p18 W=5.99u L=180.00n
MM2 ZN A1 VDD VNW p18 W=6.06u L=180.00n
.ENDS NAND2UHDV6
.SUBCKT NAND2UHDV8 A1 A2 ZN VDD VSS VNW VPW
MM3 net4 A2 VSS VPW n18 W=5.76u L=180.00n
MM1 ZN A1 net4 VPW n18 W=5.76u L=180.00n
MM0 ZN A2 VDD VNW p18 W=7.975u L=180.00n
MM2 ZN A1 VDD VNW p18 W=8.08u L=180.00n
.ENDS NAND2UHDV8
.SUBCKT NAND2XBUHDV0P4 A1 B1 ZN VDD VSS VNW VPW
MM7 net26 A1 VDD VNW p18 W=490.00n L=180.00n
MM0 ZN net26 VDD VNW p18 W=490.00n L=180.00n
MM1 ZN B1 VDD VNW p18 W=490.00n L=180.00n
MM15 net047 net26 VSS VPW n18 W=0.28u L=180.00n
MM3 net26 A1 VSS VPW n18 W=0.28u L=180.00n
MM2 ZN B1 net047 VPW n18 W=0.28u L=180.00n
.ENDS NAND2XBUHDV0P4
.SUBCKT NAND2XBUHDV0P7 A1 B1 ZN VDD VSS VNW VPW
MM15 net4 net12 VSS VPW n18 W=0.52u L=180.00n
MM2 ZN B1 net4 VPW n18 W=0.52u L=180.00n
MM3 net12 A1 VSS VPW n18 W=0.42u L=180.00n
MM1 ZN B1 VDD VNW p18 W=0.8u L=180.00n
MM0 ZN net12 VDD VNW p18 W=0.8u L=180.00n
MM7 net12 A1 VDD VNW p18 W=0.51u L=180.00n
.ENDS NAND2XBUHDV0P7
.SUBCKT NAND2XBUHDV1 A1 B1 ZN VDD VSS VNW VPW
MM15 net4 net12 VSS VPW n18 W=720.00n L=180.00n
MM2 ZN B1 net4 VPW n18 W=720.00n L=180.00n
MM3 net12 A1 VSS VPW n18 W=0.42u L=180.00n
MM1 ZN B1 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN net12 VDD VNW p18 W=1.01u L=180.00n
MM7 net12 A1 VDD VNW p18 W=0.595u L=180.00n
.ENDS NAND2XBUHDV1
.SUBCKT NAND2XBUHDV2 A1 B1 ZN VDD VSS VNW VPW
MM15 net4 net12 VSS VPW n18 W=1.44u L=180.00n
MM2 ZN B1 net4 VPW n18 W=1.44u L=180.00n
MM3 net12 A1 VSS VPW n18 W=0.59u L=180.00n
MM1 ZN B1 VDD VNW p18 W=2.02u L=180.00n
MM0 ZN net12 VDD VNW p18 W=2.02u L=180.00n
MM7 net12 A1 VDD VNW p18 W=0.97u L=180.00n
.ENDS NAND2XBUHDV2
.SUBCKT NAND2XBUHDV4 A1 B1 ZN VDD VSS VNW VPW
MM15 net4 net12 VSS VPW n18 W=2.88u L=180.00n
MM2 ZN B1 net4 VPW n18 W=2.67u L=180.00n
MM3 net12 A1 VSS VPW n18 W=0.84u L=180.00n
MM1 ZN B1 VDD VNW p18 W=4.04u L=180.00n
MM0 ZN net12 VDD VNW p18 W=3.95u L=180.00n
MM7 net12 A1 VDD VNW p18 W=1.48u L=180.00n
.ENDS NAND2XBUHDV4
.SUBCKT NAND2XBUHDV6 A1 B1 ZN VDD VSS VNW VPW
MM15 net4 net12 VSS VPW n18 W=4.32u L=180.00n
MM2 ZN B1 net4 VPW n18 W=3.9u L=180.00n
MM3 net12 A1 VSS VPW n18 W=1.44u L=180.00n
MM1 ZN B1 VDD VNW p18 W=6.06u L=180.00n
MM0 ZN net12 VDD VNW p18 W=5.88u L=180.00n
MM7 net12 A1 VDD VNW p18 W=2.02u L=180.00n
.ENDS NAND2XBUHDV6
.SUBCKT NAND2XBUHDV8 A1 B1 ZN VDD VSS VNW VPW
MM15 net4 net12 VSS VPW n18 W=5.76u L=180.00n
MM2 ZN B1 net4 VPW n18 W=5.13u L=180.00n
MM3 net12 A1 VSS VPW n18 W=1.44u L=180.00n
MM1 ZN B1 VDD VNW p18 W=8.08u L=180.00n
MM0 ZN net12 VDD VNW p18 W=7.81u L=180.00n
MM7 net12 A1 VDD VNW p18 W=2.02u L=180.00n
.ENDS NAND2XBUHDV8
.SUBCKT NAND3BBUHDV0P7 A1 A2 B ZN VDD VSS VNW VPW
MM6 net25 A2 VDD VNW p18 W=0.51u L=180.00n
MM7 net29 A1 VDD VNW p18 W=0.51u L=180.00n
MM0 ZN net25 VDD VNW p18 W=0.805u L=180.00n
MM1 ZN net29 VDD VNW p18 W=0.805u L=180.00n
MM4 ZN B VDD VNW p18 W=0.805u L=180.00n
MM8 net25 A2 VSS VPW n18 W=0.425u L=180.00n
MM3 net29 A1 VSS VPW n18 W=0.435u L=180.00n
MM2 net37 net25 net33 VPW n18 W=0.555u L=180.00n
MM15 net33 B VSS VPW n18 W=0.555u L=180.00n
MM5 ZN net29 net37 VPW n18 W=0.555u L=180.00n
.ENDS NAND3BBUHDV0P7
.SUBCKT NAND3BBUHDV1 A1 A2 B ZN VDD VSS VNW VPW
MM5 ZN net17 net9 VPW n18 W=720.00n L=180.00n
MM2 net9 net21 net13 VPW n18 W=720.00n L=180.00n
MM15 net13 B VSS VPW n18 W=720.00n L=180.00n
MM3 net17 A1 VSS VPW n18 W=0.435u L=180.00n
MM8 net21 A2 VSS VPW n18 W=0.42u L=180.00n
MM1 ZN net17 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN net21 VDD VNW p18 W=1.01u L=180.00n
MM4 ZN B VDD VNW p18 W=1.01u L=180.00n
MM7 net17 A1 VDD VNW p18 W=0.595u L=180.00n
MM6 net21 A2 VDD VNW p18 W=0.595u L=180.00n
.ENDS NAND3BBUHDV1
.SUBCKT NAND3BBUHDV2 A1 A2 B ZN VDD VSS VNW VPW
MM6 net25 A2 VDD VNW p18 W=0.595u L=180.00n
MM7 net29 A1 VDD VNW p18 W=0.97u L=180.00n
MM4 ZN B VDD VNW p18 W=2.02u L=180.00n
MM0 ZN net25 VDD VNW p18 W=1.9u L=180.00n
MM1 ZN net29 VDD VNW p18 W=1.9u L=180.00n
MM8 net25 A2 VSS VPW n18 W=0.43u L=180.00n
MM3 net29 A1 VSS VPW n18 W=0.64u L=180.00n
MM15 net33 B VSS VPW n18 W=1.44u L=180.00n
MM2 net37 net25 net33 VPW n18 W=1.44u L=180.00n
MM5 ZN net29 net37 VPW n18 W=1.44u L=180.00n
.ENDS NAND3BBUHDV2
.SUBCKT NAND3BUHDV0P7 A1 B1 B2 ZN VDD VSS VNW VPW
MM7 a1n A1 VSS VPW n18 W=0.42u L=180.00n
MM5 net9 B2 VSS VPW n18 W=0.52u L=180.00n
MM3 net13 B1 net9 VPW n18 W=0.52u L=180.00n
MM1 ZN a1n net13 VPW n18 W=0.52u L=180.00n
MM6 a1n A1 VDD VNW p18 W=0.51u L=180.00n
MM4 ZN B2 VDD VNW p18 W=0.81u L=180.00n
MM0 ZN B1 VDD VNW p18 W=0.81u L=180.00n
MM2 ZN a1n VDD VNW p18 W=0.81u L=180.00n
.ENDS NAND3BUHDV0P7
.SUBCKT NAND3BUHDV1 A1 B1 B2 ZN VDD VSS VNW VPW
MM2 ZN a1n VDD VNW p18 W=1.01u L=180.00n
MM0 ZN B1 VDD VNW p18 W=1.01u L=180.00n
MM4 ZN B2 VDD VNW p18 W=1.01u L=180.00n
MM6 a1n A1 VDD VNW p18 W=0.6u L=180.00n
MM1 ZN a1n net25 VPW n18 W=720.00n L=180.00n
MM3 net25 B1 net29 VPW n18 W=720.00n L=180.00n
MM5 net29 B2 VSS VPW n18 W=720.00n L=180.00n
MM7 a1n A1 VSS VPW n18 W=0.42u L=180.00n
.ENDS NAND3BUHDV1
.SUBCKT NAND3BUHDV2 A1 B1 B2 ZN VDD VSS VNW VPW
MM7 a1n A1 VSS VPW n18 W=0.68u L=180.00n
MM5 net9 B2 VSS VPW n18 W=1.44u L=180.00n
MM3 net13 B1 net9 VPW n18 W=1.44u L=180.00n
MM1 ZN a1n net13 VPW n18 W=1.44u L=180.00n
MM6 a1n A1 VDD VNW p18 W=0.97u L=180.00n
MM4 ZN B2 VDD VNW p18 W=1.98u L=180.00n
MM0 ZN B1 VDD VNW p18 W=1.945u L=180.00n
MM2 ZN a1n VDD VNW p18 W=1.745u L=180.00n
.ENDS NAND3BUHDV2
.SUBCKT NAND3UHDV0P4 A1 A2 A3 ZN VDD VSS VNW VPW
MM5 net5 A3 VSS VPW n18 W=0.28u L=180.00n
MM3 net9 A2 net5 VPW n18 W=0.28u L=180.00n
MM1 ZN A1 net9 VPW n18 W=0.28u L=180.00n
MM4 ZN A3 VDD VNW p18 W=0.495u L=180.00n
MM0 ZN A2 VDD VNW p18 W=0.495u L=180.00n
MM2 ZN A1 VDD VNW p18 W=0.495u L=180.00n
.ENDS NAND3UHDV0P4
.SUBCKT NAND3UHDV0P7 A1 A2 A3 ZN VDD VSS VNW VPW
MM2 ZN A1 VDD VNW p18 W=0.81u L=180.00n
MM0 ZN A2 VDD VNW p18 W=0.81u L=180.00n
MM4 ZN A3 VDD VNW p18 W=0.81u L=180.00n
MM1 ZN A1 net21 VPW n18 W=0.61u L=180.00n
MM3 net21 A2 net25 VPW n18 W=0.61u L=180.00n
MM5 net25 A3 VSS VPW n18 W=0.61u L=180.00n
.ENDS NAND3UHDV0P7
.SUBCKT NAND3UHDV1 A1 A2 A3 ZN VDD VSS VNW VPW
MM2 ZN A1 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN A2 VDD VNW p18 W=1.01u L=180.00n
MM4 ZN A3 VDD VNW p18 W=1.01u L=180.00n
MM1 ZN A1 net21 VPW n18 W=720.00n L=180.00n
MM3 net21 A2 net25 VPW n18 W=720.00n L=180.00n
MM5 net25 A3 VSS VPW n18 W=720.00n L=180.00n
.ENDS NAND3UHDV1
.SUBCKT NAND3UHDV2 A1 A2 A3 ZN VDD VSS VNW VPW
MM2 ZN A1 VDD VNW p18 W=1.9u L=180.00n
MM0 ZN A2 VDD VNW p18 W=1.9u L=180.00n
MM4 ZN A3 VDD VNW p18 W=2.02u L=180.00n
MM1 ZN A1 net21 VPW n18 W=1.44u L=180.00n
MM3 net21 A2 net25 VPW n18 W=1.44u L=180.00n
MM5 net25 A3 VSS VPW n18 W=1.44u L=180.00n
.ENDS NAND3UHDV2
.SUBCKT NAND4BUHDV0P7 A1 B1 B2 B3 ZN VDD VSS VNW VPW
MM7 ZN net26 VDD VNW p18 W=0.78u L=180.00n
MM8 net26 A1 VDD VNW p18 W=0.49u L=180.00n
MM2 ZN B1 VDD VNW p18 W=0.78u L=180.00n
MM0 ZN B2 VDD VNW p18 W=0.78u L=180.00n
MM4 ZN B3 VDD VNW p18 W=0.78u L=180.00n
MM9 net26 A1 VSS VPW n18 W=0.49u L=180.00n
MM6 ZN net26 net30 VPW n18 W=0.61u L=180.00n
MM1 net30 B1 net34 VPW n18 W=0.61u L=180.00n
MM3 net34 B2 net38 VPW n18 W=0.61u L=180.00n
MM5 net38 B3 VSS VPW n18 W=0.61u L=180.00n
.ENDS NAND4BUHDV0P7
.SUBCKT NAND4BUHDV1 A1 B1 B2 B3 ZN VDD VSS VNW VPW
MM6 ZN net22 net18 VPW n18 W=720.00n L=180.00n
MM5 net10 B3 VSS VPW n18 W=720.00n L=180.00n
MM3 net14 B2 net10 VPW n18 W=720.00n L=180.00n
MM1 net18 B1 net14 VPW n18 W=720.00n L=180.00n
MM9 net22 A1 VSS VPW n18 W=440.00n L=180.00n
MM4 ZN B3 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN B2 VDD VNW p18 W=1.01u L=180.00n
MM2 ZN B1 VDD VNW p18 W=1.01u L=180.00n
MM7 ZN net22 VDD VNW p18 W=1.01u L=180.00n
MM8 net22 A1 VDD VNW p18 W=580.0n L=180.00n
.ENDS NAND4BUHDV1
.SUBCKT NAND4BUHDV2 A1 B1 B2 B3 ZN VDD VSS VNW VPW
MM6 ZN net22 net18 VPW n18 W=1.44u L=180.00n
MM5 net10 B3 VSS VPW n18 W=1220.00n L=180.00n
MM3 net14 B2 net10 VPW n18 W=1.44u L=180.00n
MM1 net18 B1 net14 VPW n18 W=1.44u L=180.00n
MM9 net22 A1 VSS VPW n18 W=0.68u L=180.00n
MM4 ZN B3 VDD VNW p18 W=2.02u L=180.00n
MM0 ZN B2 VDD VNW p18 W=2.02u L=180.00n
MM2 ZN B1 VDD VNW p18 W=1.96u L=180.00n
MM7 ZN net22 VDD VNW p18 W=1.96u L=180.00n
MM8 net22 A1 VDD VNW p18 W=950.0n L=180.00n
.ENDS NAND4BUHDV2
.SUBCKT NAND4UHDV0P7 A1 A2 A3 A4 ZN VDD VSS VNW VPW
MM5 net6 A4 VSS VPW n18 W=560.00n L=180.00n
MM3 net10 A3 net6 VPW n18 W=560.00n L=180.00n
MM1 net14 A2 net10 VPW n18 W=560.00n L=180.00n
MM6 ZN A1 net14 VPW n18 W=560.00n L=180.00n
MM4 ZN A4 VDD VNW p18 W=0.475u L=180.00n
MM0 ZN A3 VDD VNW p18 W=0.475u L=180.00n
MM2 ZN A2 VDD VNW p18 W=0.475u L=180.00n
MM7 ZN A1 VDD VNW p18 W=0.475u L=180.00n
.ENDS NAND4UHDV0P7
.SUBCKT NAND4UHDV1 A1 A2 A3 A4 ZN VDD VSS VNW VPW
MM7 ZN A1 VDD VNW p18 W=1.01u L=180.00n
MM2 ZN A2 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN A3 VDD VNW p18 W=1.01u L=180.00n
MM4 ZN A4 VDD VNW p18 W=1.01u L=180.00n
MM6 ZN A1 net26 VPW n18 W=720.00n L=180.00n
MM1 net26 A2 net30 VPW n18 W=720.00n L=180.00n
MM3 net30 A3 net34 VPW n18 W=720.00n L=180.00n
MM5 net34 A4 VSS VPW n18 W=720.00n L=180.00n
.ENDS NAND4UHDV1
.SUBCKT NAND4UHDV2 A1 A2 A3 A4 ZN VDD VSS VNW VPW
MM5 net6 A4 VSS VPW n18 W=1.44u L=180.00n
MM3 net10 A3 net6 VPW n18 W=1.44u L=180.00n
MM1 net14 A2 net10 VPW n18 W=1.44u L=180.00n
MM6 ZN A1 net14 VPW n18 W=1.44u L=180.00n
MM4 ZN A4 VDD VNW p18 W=2.02u L=180.00n
MM0 ZN A3 VDD VNW p18 W=2.02u L=180.00n
MM2 ZN A2 VDD VNW p18 W=1.9u L=180.00n
MM7 ZN A1 VDD VNW p18 W=1.9u L=180.00n
.ENDS NAND4UHDV2
.SUBCKT NAND4XXBBUHDV0P7 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM5 net032 A1 VSS VPW n18 W=0.475u L=180.00n
MM6 ZN B1 net22 VPW n18 W=0.605u L=180.00n
MM3 net18 net032 VSS VPW n18 W=0.605u L=180.00n
MM1 net22 B2 net18 VPW n18 W=0.605u L=180.00n
MM9 net032 A2 VSS VPW n18 W=0.475u L=180.00n
MM4 net33 A1 VDD VNW p18 W=0.515u L=180.00n
MM0 ZN B2 VDD VNW p18 W=0.805u L=180.00n
MM2 ZN B1 VDD VNW p18 W=0.805u L=180.00n
MM7 ZN net032 VDD VNW p18 W=0.805u L=180.00n
MM8 net032 A2 net33 VNW p18 W=0.515u L=180.00n
.ENDS NAND4XXBBUHDV0P7
.SUBCKT NAND4XXBBUHDV1 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM7 ZN net30 VDD VNW p18 W=1.01u L=180.00n
MM2 ZN B1 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN B2 VDD VNW p18 W=1.01u L=180.00n
MM8 net30 A2 net21 VNW p18 W=0.595u L=180.00n
MM4 net21 A1 VDD VNW p18 W=0.595u L=180.00n
MM9 net30 A2 VSS VPW n18 W=0.475u L=180.00n
MM5 net30 A1 VSS VPW n18 W=0.475u L=180.00n
MM1 net34 B2 net38 VPW n18 W=720.00n L=180.00n
MM3 net38 net30 VSS VPW n18 W=720.00n L=180.00n
MM6 ZN B1 net34 VPW n18 W=720.00n L=180.00n
.ENDS NAND4XXBBUHDV1
.SUBCKT NAND4XXBBUHDV2 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM7 ZN net30 VDD VNW p18 W=2.02u L=180.00n
MM2 ZN B1 VDD VNW p18 W=1.9u L=180.00n
MM0 ZN B2 VDD VNW p18 W=2.02u L=180.00n
MM8 net30 A2 net21 VNW p18 W=0.97u L=180.00n
MM4 net21 A1 VDD VNW p18 W=0.97u L=180.00n
MM9 net30 A2 VSS VPW n18 W=0.7u L=180.00n
MM5 net30 A1 VSS VPW n18 W=0.7u L=180.00n
MM1 net34 B2 net38 VPW n18 W=1.44u L=180.00n
MM3 net38 net30 VSS VPW n18 W=1.44u L=180.00n
MM6 ZN B1 net34 VPW n18 W=1.44u L=180.00n
.ENDS NAND4XXBBUHDV2
.SUBCKT NAND4XXBBUHDV3 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM7 ZN net30 VDD VNW p18 W=3.03u L=180.00n
MM2 ZN B1 VDD VNW p18 W=2.72u L=180.00n
MM0 ZN B2 VDD VNW p18 W=2.655u L=180.00n
MM8 net30 A2 net21 VNW p18 W=1.01u L=180.00n
MM4 net21 A1 VDD VNW p18 W=1.01u L=180.00n
MM9 net30 A2 VSS VPW n18 W=0.72u L=180.00n
MM5 net30 A1 VSS VPW n18 W=0.72u L=180.00n
MM1 net34 B2 net38 VPW n18 W=2.16u L=180.00n
MM3 net38 net30 VSS VPW n18 W=2.16u L=180.00n
MM6 ZN B1 net34 VPW n18 W=2.16u L=180.00n
.ENDS NAND4XXBBUHDV3
.SUBCKT NDQUHDV0P7 CKN D Q VDD VSS VNW VPW
MM6 net88 c net55 VNW p18 W=0.59u L=180.00n
MM11 net56 net55 VDD VNW p18 W=0.59u L=180.00n
MM12 net19 net56 VDD VNW p18 W=0.59u L=180.00n
MM14 net55 cn net19 VNW p18 W=0.59u L=180.00n
MM26 net68 c net79 VNW p18 W=0.89u L=180.00n
MM25 Q net92 VDD VNW p18 W=0.8u L=180.00n
MM17 net56 cn net79 VNW p18 W=590.00n L=180.00n
MM1 c CKN VDD VNW p18 W=420.00n L=180.00n
MM3 cn c VDD VNW p18 W=250.00n L=180.00n
MM5 net88 D VDD VNW p18 W=0.59u L=180.00n
MM23 net92 net79 VDD VNW p18 W=1.01u L=180.00n
MM22 net68 net92 VDD VNW p18 W=0.95u L=180.00n
MM9 net88 cn net55 VPW n18 W=0.6u L=180.00n
MM10 net56 net55 VSS VPW n18 W=0.34u L=180.00n
MM13 net55 c net64 VPW n18 W=0.73u L=180.00n
MM15 net64 net56 VSS VPW n18 W=0.34u L=180.00n
MM31 net68 cn net79 VPW n18 W=430.00n L=180.00n
MM24 Q net92 VSS VPW n18 W=0.57u L=180.00n
MM16 net56 c net79 VPW n18 W=430.00n L=180.00n
MM0 c CKN VSS VPW n18 W=360.00n L=180.00n
MM2 cn c VSS VPW n18 W=420.00n L=180.00n
MM4 net88 D VSS VPW n18 W=0.34u L=180.00n
MM20 net92 net79 VSS VPW n18 W=590.00n L=180.00n
MM18 net68 net92 VSS VPW n18 W=430.00n L=180.00n
.ENDS NDQUHDV0P7
.SUBCKT NDQUHDV1 CKN D Q VDD VSS VNW VPW
MM18 net32 net8 VSS VPW n18 W=430.00n L=180.00n
MM20 net8 net27 VSS VPW n18 W=590.00n L=180.00n
MM4 net12 D VSS VPW n18 W=0.34u L=180.00n
MM2 cn c VSS VPW n18 W=420.00n L=180.00n
MM0 c CKN VSS VPW n18 W=250.00n L=180.00n
MM16 net44 c net27 VPW n18 W=430.00n L=180.00n
MM24 Q net8 VSS VPW n18 W=720.00n L=180.00n
MM31 net32 cn net27 VPW n18 W=430.00n L=180.00n
MM15 net36 net44 VSS VPW n18 W=0.34u L=180.00n
MM13 net51 c net36 VPW n18 W=0.73u L=180.00n
MM10 net44 net51 VSS VPW n18 W=0.34u L=180.00n
MM9 net12 cn net51 VPW n18 W=0.6u L=180.00n
MM22 net32 net8 VDD VNW p18 W=0.95u L=180.00n
MM23 net8 net27 VDD VNW p18 W=1.01u L=180.00n
MM5 net12 D VDD VNW p18 W=0.59u L=180.00n
MM3 cn c VDD VNW p18 W=250.00n L=180.00n
MM1 c CKN VDD VNW p18 W=420.00n L=180.00n
MM17 net44 cn net27 VNW p18 W=590.00n L=180.00n
MM25 Q net8 VDD VNW p18 W=1.01u L=180.00n
MM26 net32 c net27 VNW p18 W=0.89u L=180.00n
MM14 net51 cn net87 VNW p18 W=0.59u L=180.00n
MM11 net44 net51 VDD VNW p18 W=0.59u L=180.00n
MM6 net12 c net51 VNW p18 W=0.59u L=180.00n
MM12 net87 net44 VDD VNW p18 W=0.59u L=180.00n
.ENDS NDQUHDV1
.SUBCKT NDQUHDV2 CKN D Q VDD VSS VNW VPW
MM18 net32 net8 VSS VPW n18 W=0.53u L=180.00n
MM20 net8 net27 VSS VPW n18 W=0.53u L=180.00n
MM4 net12 D VSS VPW n18 W=0.34u L=180.00n
MM2 cn c VSS VPW n18 W=420.00n L=180.00n
MM0 c CKN VSS VPW n18 W=250.00n L=180.00n
MM16 net44 c net27 VPW n18 W=0.53u L=180.00n
MM24 Q net8 VSS VPW n18 W=1.44u L=180.00n
MM31 net32 cn net27 VPW n18 W=0.53u L=180.00n
MM15 net36 net44 VSS VPW n18 W=0.34u L=180.00n
MM13 net51 c net36 VPW n18 W=0.73u L=180.00n
MM10 net44 net51 VSS VPW n18 W=0.34u L=180.00n
MM9 net12 cn net51 VPW n18 W=0.6u L=180.00n
MM22 net32 net8 VDD VNW p18 W=0.95u L=180.00n
MM23 net8 net27 VDD VNW p18 W=1.01u L=180.00n
MM5 net12 D VDD VNW p18 W=0.59u L=180.00n
MM3 cn c VDD VNW p18 W=250.00n L=180.00n
MM1 c CKN VDD VNW p18 W=420.00n L=180.00n
MM17 net44 cn net27 VNW p18 W=590.00n L=180.00n
MM25 Q net8 VDD VNW p18 W=2.02u L=180.00n
MM26 net32 c net27 VNW p18 W=0.89u L=180.00n
MM14 net51 cn net87 VNW p18 W=0.59u L=180.00n
MM11 net44 net51 VDD VNW p18 W=0.59u L=180.00n
MM6 net12 c net51 VNW p18 W=0.59u L=180.00n
MM12 net87 net44 VDD VNW p18 W=0.59u L=180.00n
.ENDS NDQUHDV2
.SUBCKT NDQUHDV3 CKN D Q VDD VSS VNW VPW
MM12 net19 net56 VDD VNW p18 W=0.59u L=180.00n
MM6 net88 c net55 VNW p18 W=0.59u L=180.00n
MM11 net56 net55 VDD VNW p18 W=0.59u L=180.00n
MM14 net55 cn net19 VNW p18 W=0.59u L=180.00n
MM26 net68 c net79 VNW p18 W=0.89u L=180.00n
MM25 Q net92 VDD VNW p18 W=3.03u L=180.00n
MM17 net56 cn net79 VNW p18 W=590.00n L=180.00n
MM1 c CKN VDD VNW p18 W=420.00n L=180.00n
MM3 cn c VDD VNW p18 W=250.00n L=180.00n
MM5 net88 D VDD VNW p18 W=0.59u L=180.00n
MM23 net92 net79 VDD VNW p18 W=1.01u L=180.00n
MM22 net68 net92 VDD VNW p18 W=0.95u L=180.00n
MM9 net88 cn net55 VPW n18 W=0.6u L=180.00n
MM10 net56 net55 VSS VPW n18 W=0.34u L=180.00n
MM13 net55 c net64 VPW n18 W=0.73u L=180.00n
MM15 net64 net56 VSS VPW n18 W=0.34u L=180.00n
MM31 net68 cn net79 VPW n18 W=0.53u L=180.00n
MM24 Q net92 VSS VPW n18 W=2.16u L=180.00n
MM16 net56 c net79 VPW n18 W=0.53u L=180.00n
MM0 c CKN VSS VPW n18 W=250.00n L=180.00n
MM2 cn c VSS VPW n18 W=420.00n L=180.00n
MM4 net88 D VSS VPW n18 W=0.34u L=180.00n
MM20 net92 net79 VSS VPW n18 W=0.53u L=180.00n
MM18 net68 net92 VSS VPW n18 W=0.53u L=180.00n
.ENDS NDQUHDV3
.SUBCKT NDSRNQUHDV1 CKN D Q RDN SDN VDD VSS VNW VPW
MM29 net108 c net61 VNW p18 W=0.42u L=180.00n
MM30 net101 SDN VDD VNW p18 W=0.37u L=180.00n
MM32 net108 cn net88 VNW p18 W=0.42u L=180.00n
MM21 net88 net101 VDD VNW p18 W=0.42u L=180.00n
MM20 net88 RDN VDD VNW p18 W=0.42u L=180.00n
MM14 net101 cn net100 VNW p18 W=0.425u L=180.00n
MM10 net101 net108 VDD VNW p18 W=0.42u L=180.00n
MM6 cn c VDD VNW p18 W=250.00n L=180.00n
MM2 c CKN VDD VNW p18 W=420.00n L=180.00n
MM0 net61 D VDD VNW p18 W=0.42u L=180.00n
MM16 net112 RDN VDD VNW p18 W=0.35u L=180.00n
MM17 net112 net100 VDD VNW p18 W=0.35u L=180.00n
MM5 Q net112 VDD VNW p18 W=1.01u L=180.00n
MM34 net0204 net112 VDD VNW p18 W=0.42u L=180.00n
MM35 net0204 SDN VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net0204 VNW p18 W=0.425u L=180.00n
MM37 net100 cn net0264 VPW n18 W=0.42u L=180.00n
MM38 net0264 SDN net0260 VPW n18 W=0.42u L=180.00n
MM33 net108 c net0292 VPW n18 W=0.445u L=180.00n
MM31 net0276 net108 VSS VPW n18 W=0.49u L=180.00n
MM28 net108 cn net0320 VPW n18 W=0.445u L=180.00n
MM39 net0260 net112 VSS VPW n18 W=0.42u L=180.00n
MM1 net0320 D VSS VPW n18 W=0.445u L=180.00n
MM7 cn c VSS VPW n18 W=420.00n L=180.00n
MM3 c CKN VSS VPW n18 W=250.00n L=180.00n
MM19 net112 net100 net77 VPW n18 W=0.53u L=180.00n
MM18 net77 RDN VSS VPW n18 W=0.53u L=180.00n
MM23 net0292 RDN net93 VPW n18 W=0.445u L=180.00n
MM22 net93 net101 VSS VPW n18 W=0.445u L=180.00n
MM15 net101 c net100 VPW n18 W=0.42u L=180.00n
MM12 net101 SDN net0276 VPW n18 W=0.49u L=180.00n
MM4 Q net112 VSS VPW n18 W=0.72u L=180.00n
.ENDS NDSRNQUHDV1
.SUBCKT NDSRNQUHDV2 CKN D Q RDN SDN VDD VSS VNW VPW
MM29 net108 c net61 VNW p18 W=0.42u L=180.00n
MM30 net101 SDN VDD VNW p18 W=0.37u L=180.00n
MM32 net108 cn net88 VNW p18 W=0.42u L=180.00n
MM21 net88 net101 VDD VNW p18 W=0.42u L=180.00n
MM20 net88 RDN VDD VNW p18 W=0.42u L=180.00n
MM14 net101 cn net100 VNW p18 W=0.425u L=180.00n
MM10 net101 net108 VDD VNW p18 W=0.42u L=180.00n
MM6 cn c VDD VNW p18 W=250.00n L=180.00n
MM2 c CKN VDD VNW p18 W=420.00n L=180.00n
MM0 net61 D VDD VNW p18 W=0.42u L=180.00n
MM16 net112 RDN VDD VNW p18 W=0.35u L=180.00n
MM17 net112 net100 VDD VNW p18 W=0.43u L=180.00n
MM5 Q net112 VDD VNW p18 W=2.02u L=180.00n
MM34 net0204 net112 VDD VNW p18 W=0.42u L=180.00n
MM35 net0204 SDN VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net0204 VNW p18 W=0.425u L=180.00n
MM37 net100 cn net0264 VPW n18 W=0.42u L=180.00n
MM38 net0264 SDN net0260 VPW n18 W=0.42u L=180.00n
MM33 net108 c net0292 VPW n18 W=0.445u L=180.00n
MM31 net0276 net108 VSS VPW n18 W=0.49u L=180.00n
MM28 net108 cn net0320 VPW n18 W=0.445u L=180.00n
MM39 net0260 net112 VSS VPW n18 W=0.42u L=180.00n
MM1 net0320 D VSS VPW n18 W=0.445u L=180.00n
MM7 cn c VSS VPW n18 W=420.00n L=180.00n
MM3 c CKN VSS VPW n18 W=250.00n L=180.00n
MM19 net112 net100 net77 VPW n18 W=0.53u L=180.00n
MM18 net77 RDN VSS VPW n18 W=0.53u L=180.00n
MM23 net0292 RDN net93 VPW n18 W=0.445u L=180.00n
MM22 net93 net101 VSS VPW n18 W=0.445u L=180.00n
MM15 net101 c net100 VPW n18 W=0.42u L=180.00n
MM12 net101 SDN net0276 VPW n18 W=0.49u L=180.00n
MM4 Q net112 VSS VPW n18 W=1.44u L=180.00n
.ENDS NDSRNQUHDV2
.SUBCKT NOR2UHDV0P4 A1 A2 ZN VDD VSS VNW VPW
MM5 ZN A2 VSS VPW n18 W=0.28u L=180.00n
MM9 ZN A1 VSS VPW n18 W=0.28u L=180.00n
MM4 net19 A2 VDD VNW p18 W=490.0n L=180.00n
MM8 ZN A1 net19 VNW p18 W=490.0n L=180.00n
.ENDS NOR2UHDV0P4
.SUBCKT NOR2UHDV0P7 A1 A2 ZN VDD VSS VNW VPW
MM8 ZN A1 net7 VNW p18 W=790.0n L=180.00n
MM4 net7 A2 VDD VNW p18 W=790.0n L=180.00n
MM9 ZN A1 VSS VPW n18 W=560.00n L=180.00n
MM5 ZN A2 VSS VPW n18 W=560.00n L=180.00n
.ENDS NOR2UHDV0P7
.SUBCKT NOR2UHDV1 A1 A2 ZN VDD VSS VNW VPW
MM8 ZN A1 net7 VNW p18 W=1.01u L=180.00n
MM4 net7 A2 VDD VNW p18 W=1.01u L=180.00n
MM9 ZN A1 VSS VPW n18 W=720.00n L=180.00n
MM5 ZN A2 VSS VPW n18 W=720.00n L=180.00n
.ENDS NOR2UHDV1
.SUBCKT NOR2UHDV2 A1 A2 ZN VDD VSS VNW VPW
MM8 ZN A1 net7 VNW p18 W=2.02u L=180.00n
MM4 net7 A2 VDD VNW p18 W=2.02u L=180.00n
MM9 ZN A1 VSS VPW n18 W=1.44u L=180.00n
MM5 ZN A2 VSS VPW n18 W=1.44u L=180.00n
.ENDS NOR2UHDV2
.SUBCKT NOR2UHDV3 A1 A2 ZN VDD VSS VNW VPW
MM8 ZN A1 net7 VNW p18 W=3.03u L=180.00n
MM4 net7 A2 VDD VNW p18 W=2.995u L=180.00n
MM9 ZN A1 VSS VPW n18 W=2.14u L=180.00n
MM5 ZN A2 VSS VPW n18 W=2.14u L=180.00n
.ENDS NOR2UHDV3
.SUBCKT NOR2UHDV4 A1 A2 ZN VDD VSS VNW VPW
MM8 ZN A1 net7 VNW p18 W=4.04u L=180.00n
MM4 net7 A2 VDD VNW p18 W=3.8u L=180.00n
MM9 ZN A1 VSS VPW n18 W=2.88u L=180.00n
MM5 ZN A2 VSS VPW n18 W=2.88u L=180.00n
.ENDS NOR2UHDV4
.SUBCKT NOR2UHDV6 A1 A2 ZN VDD VSS VNW VPW
MM8 ZN A1 net7 VNW p18 W=6.06u L=180.00n
MM4 net7 A2 VDD VNW p18 W=5.785u L=180.00n
MM9 ZN A1 VSS VPW n18 W=4.32u L=180.00n
MM5 ZN A2 VSS VPW n18 W=4.32u L=180.00n
.ENDS NOR2UHDV6
.SUBCKT NOR2UHDV8 A1 A2 ZN VDD VSS VNW VPW
MM8 ZN A1 net7 VNW p18 W=8.08u L=180.00n
MM4 net7 A2 VDD VNW p18 W=7.77u L=180.00n
MM9 ZN A1 VSS VPW n18 W=5.76u L=180.00n
MM5 ZN A2 VSS VPW n18 W=5.76u L=180.00n
.ENDS NOR2UHDV8
.SUBCKT NOR2XBUHDV0P4 A1 B1 ZN VDD VSS VNW VPW
MM4 ZN B1 net11 VNW p18 W=490.0n L=180.00n
MM2 net11 net24 VDD VNW p18 W=490.0n L=180.00n
MM1 net24 A1 VDD VNW p18 W=490.0n L=180.00n
MM5 ZN B1 VSS VPW n18 W=0.28u L=180.00n
MM3 ZN net24 VSS VPW n18 W=0.28u L=180.00n
MM0 net24 A1 VSS VPW n18 W=0.28u L=180.00n
.ENDS NOR2XBUHDV0P4
.SUBCKT NOR2XBUHDV0P7 A1 B1 ZN VDD VSS VNW VPW
MM0 net4 A1 VSS VPW n18 W=430.00n L=180.00n
MM3 ZN net4 VSS VPW n18 W=560.00n L=180.00n
MM5 ZN B1 VSS VPW n18 W=560.00n L=180.00n
MM1 net4 A1 VDD VNW p18 W=500.0n L=180.00n
MM4 ZN B1 net23 VNW p18 W=790.0n L=180.00n
MM2 net23 net4 VDD VNW p18 W=790.0n L=180.00n
.ENDS NOR2XBUHDV0P7
.SUBCKT NOR2XBUHDV1 A1 B1 ZN VDD VSS VNW VPW
MM2 net11 net24 VDD VNW p18 W=1.01u L=180.00n
MM4 ZN B1 net11 VNW p18 W=1.01u L=180.00n
MM1 net24 A1 VDD VNW p18 W=580.0n L=180.00n
MM5 ZN B1 VSS VPW n18 W=720.00n L=180.00n
MM3 ZN net24 VSS VPW n18 W=720.00n L=180.00n
MM0 net24 A1 VSS VPW n18 W=430.00n L=180.00n
.ENDS NOR2XBUHDV1
.SUBCKT NOR2XBUHDV2 A1 B1 ZN VDD VSS VNW VPW
MM0 net4 A1 VSS VPW n18 W=690.00n L=180.00n
MM3 ZN net4 VSS VPW n18 W=1.44u L=180.00n
MM5 ZN B1 VSS VPW n18 W=1.44u L=180.00n
MM1 net4 A1 VDD VNW p18 W=950.0n L=180.00n
MM4 ZN B1 net23 VNW p18 W=2.02u L=180.00n
MM2 net23 net4 VDD VNW p18 W=2.02u L=180.00n
.ENDS NOR2XBUHDV2
.SUBCKT NOR2XBUHDV3 A1 B1 ZN VDD VSS VNW VPW
MM0 net4 A1 VSS VPW n18 W=720.00n L=180.00n
MM3 ZN net4 VSS VPW n18 W=2.16u L=180.00n
MM5 ZN B1 VSS VPW n18 W=2.16u L=180.00n
MM1 net4 A1 VDD VNW p18 W=1.01u L=180.00n
MM4 ZN B1 net23 VNW p18 W=3.03u L=180.00n
MM2 net23 net4 VDD VNW p18 W=2.85u L=180.00n
.ENDS NOR2XBUHDV3
.SUBCKT NOR2XBUHDV4 A1 B1 ZN VDD VSS VNW VPW
MM0 net4 A1 VSS VPW n18 W=1060.00n L=180.00n
MM3 ZN net4 VSS VPW n18 W=2.88u L=180.00n
MM5 ZN B1 VSS VPW n18 W=2.88u L=180.00n
MM1 net4 A1 VDD VNW p18 W=1.49u L=180.00n
MM4 ZN B1 net23 VNW p18 W=4.04u L=180.00n
MM2 net23 net4 VDD VNW p18 W=4.04u L=180.00n
.ENDS NOR2XBUHDV4
.SUBCKT NOR2XBUHDV6 A1 B1 ZN VDD VSS VNW VPW
MM0 net4 A1 VSS VPW n18 W=1.44u L=180.00n
MM3 ZN net4 VSS VPW n18 W=4.32u L=180.00n
MM5 ZN B1 VSS VPW n18 W=4.32u L=180.00n
MM1 net4 A1 VDD VNW p18 W=2.02u L=180.00n
MM4 ZN B1 net23 VNW p18 W=6.06u L=180.00n
MM2 net23 net4 VDD VNW p18 W=6.06u L=180.00n
.ENDS NOR2XBUHDV6
.SUBCKT NOR2XBUHDV8 A1 B1 ZN VDD VSS VNW VPW
MM0 net4 A1 VSS VPW n18 W=2.16u L=180.00n
MM3 ZN net4 VSS VPW n18 W=5.76u L=180.00n
MM5 ZN B1 VSS VPW n18 W=5.76u L=180.00n
MM1 net4 A1 VDD VNW p18 W=3.03u L=180.00n
MM4 ZN B1 net23 VNW p18 W=8.08u L=180.00n
MM2 net23 net4 VDD VNW p18 W=8.08u L=180.00n
.ENDS NOR2XBUHDV8
.SUBCKT NOR3BUHDV0P7 A1 B1 B2 ZN VDD VSS VNW VPW
MM8 net20 B1 net12 VNW p18 W=790.0n L=180.00n
MM4 net12 B2 VDD VNW p18 W=790.0n L=180.00n
MM0 ZN net21 net20 VNW p18 W=790.0n L=180.00n
MM2 net21 A1 VDD VNW p18 W=500.0n L=180.00n
MM3 net21 A1 VSS VPW n18 W=430.00n L=180.00n
MM1 ZN net21 VSS VPW n18 W=560.00n L=180.00n
MM9 ZN B1 VSS VPW n18 W=560.00n L=180.00n
MM5 ZN B2 VSS VPW n18 W=560.00n L=180.00n
.ENDS NOR3BUHDV0P7
.SUBCKT NOR3BUHDV1 A1 B1 B2 ZN VDD VSS VNW VPW
MM9 ZN B1 VSS VPW n18 W=720.00n L=180.00n
MM5 ZN B2 VSS VPW n18 W=720.00n L=180.00n
MM1 ZN net17 VSS VPW n18 W=720.00n L=180.00n
MM3 net17 A1 VSS VPW n18 W=430.00n L=180.00n
MM0 ZN net17 net24 VNW p18 W=1.01u L=180.00n
MM4 net32 B2 VDD VNW p18 W=1.01u L=180.00n
MM8 net24 B1 net32 VNW p18 W=1.01u L=180.00n
MM2 net17 A1 VDD VNW p18 W=580.0n L=180.00n
.ENDS NOR3BUHDV1
.SUBCKT NOR3BUHDV2 A1 B1 B2 ZN VDD VSS VNW VPW
MM2 net21 A1 VDD VNW p18 W=950.0n L=180.00n
MM8 net20 B1 net12 VNW p18 W=1.985u L=180.00n
MM4 net12 B2 VDD VNW p18 W=1.985u L=180.00n
MM0 ZN net21 net20 VNW p18 W=2.02u L=180.00n
MM3 net21 A1 VSS VPW n18 W=630.00n L=180.00n
MM1 ZN net21 VSS VPW n18 W=1.44u L=180.00n
MM5 ZN B2 VSS VPW n18 W=1.44u L=180.00n
MM9 ZN B1 VSS VPW n18 W=1.44u L=180.00n
.ENDS NOR3BUHDV2
.SUBCKT NOR3BUHDV3 A1 B1 B2 ZN VDD VSS VNW VPW
MM9 ZN B1 VSS VPW n18 W=2.16u L=180.00n
MM5 ZN B2 VSS VPW n18 W=2.16u L=180.00n
MM1 ZN net17 VSS VPW n18 W=2.16u L=180.00n
MM3 net17 A1 VSS VPW n18 W=720.00n L=180.00n
MM0 ZN net17 net24 VNW p18 W=3.03u L=180.00n
MM4 net32 B2 VDD VNW p18 W=3.03u L=180.00n
MM8 net24 B1 net32 VNW p18 W=3.03u L=180.00n
MM2 net17 A1 VDD VNW p18 W=1.01u L=180.00n
.ENDS NOR3BUHDV3
.SUBCKT NOR3BUHDV4 A1 B1 B2 ZN VDD VSS VNW VPW
MM2 net21 A1 VDD VNW p18 W=1.33u L=180.00n
MM8 net20 B1 net12 VNW p18 W=4.04u L=180.00n
MM4 net12 B2 VDD VNW p18 W=4.04u L=180.00n
MM0 ZN net21 net20 VNW p18 W=4.04u L=180.00n
MM3 net21 A1 VSS VPW n18 W=1060.00n L=180.00n
MM1 ZN net21 VSS VPW n18 W=2.88u L=180.00n
MM5 ZN B2 VSS VPW n18 W=2.88u L=180.00n
MM9 ZN B1 VSS VPW n18 W=2.88u L=180.00n
.ENDS NOR3BUHDV4
.SUBCKT NOR3UHDV0P4 A1 A2 A3 ZN VDD VSS VNW VPW
MM0 ZN A1 net16 VNW p18 W=490.0n L=180.00n
MM8 net16 A2 net8 VNW p18 W=490.0n L=180.00n
MM4 net8 A3 VDD VNW p18 W=490.0n L=180.00n
MM1 ZN A1 VSS VPW n18 W=0.28u L=180.00n
MM9 ZN A2 VSS VPW n18 W=0.28u L=180.00n
MM5 ZN A3 VSS VPW n18 W=0.28u L=180.00n
.ENDS NOR3UHDV0P4
.SUBCKT NOR3UHDV0P7 A1 A2 A3 ZN VDD VSS VNW VPW
MM5 ZN A3 VSS VPW n18 W=0.465u L=180.00n
MM9 ZN A2 VSS VPW n18 W=0.465u L=180.00n
MM1 ZN A1 VSS VPW n18 W=0.465u L=180.00n
MM0 ZN A1 net20 VNW p18 W=790.0n L=180.00n
MM4 net28 A3 VDD VNW p18 W=790.0n L=180.00n
MM8 net20 A2 net28 VNW p18 W=790.0n L=180.00n
.ENDS NOR3UHDV0P7
.SUBCKT NOR3UHDV1 A1 A2 A3 ZN VDD VSS VNW VPW
MM5 ZN A3 VSS VPW n18 W=720.00n L=180.00n
MM9 ZN A2 VSS VPW n18 W=720.00n L=180.00n
MM1 ZN A1 VSS VPW n18 W=720.00n L=180.00n
MM0 ZN A1 net20 VNW p18 W=1.01u L=180.00n
MM4 net28 A3 VDD VNW p18 W=1.01u L=180.00n
MM8 net20 A2 net28 VNW p18 W=1.01u L=180.00n
.ENDS NOR3UHDV1
.SUBCKT NOR3UHDV2 A1 A2 A3 ZN VDD VSS VNW VPW
MM5 ZN A3 VSS VPW n18 W=1.44u L=180.00n
MM9 ZN A2 VSS VPW n18 W=1.44u L=180.00n
MM1 ZN A1 VSS VPW n18 W=1.44u L=180.00n
MM0 ZN A1 net20 VNW p18 W=2.02u L=180.00n
MM4 net28 A3 VDD VNW p18 W=2.02u L=180.00n
MM8 net20 A2 net28 VNW p18 W=1.985u L=180.00n
.ENDS NOR3UHDV2
.SUBCKT NOR3UHDV3 A1 A2 A3 ZN VDD VSS VNW VPW
MM5 ZN A3 VSS VPW n18 W=2.16u L=180.00n
MM9 ZN A2 VSS VPW n18 W=2.16u L=180.00n
MM1 ZN A1 VSS VPW n18 W=2.16u L=180.00n
MM0 ZN A1 net20 VNW p18 W=3.03u L=180.00n
MM4 net28 A3 VDD VNW p18 W=3.03u L=180.00n
MM8 net20 A2 net28 VNW p18 W=2.99u L=180.00n
.ENDS NOR3UHDV3
.SUBCKT NOR3UHDV4 A1 A2 A3 ZN VDD VSS VNW VPW
MM5 ZN A3 VSS VPW n18 W=2.88u L=180.00n
MM9 ZN A2 VSS VPW n18 W=2.88u L=180.00n
MM1 ZN A1 VSS VPW n18 W=2.88u L=180.00n
MM0 ZN A1 net20 VNW p18 W=4.04u L=180.00n
MM4 net28 A3 VDD VNW p18 W=4.04u L=180.00n
MM8 net20 A2 net28 VNW p18 W=4u L=180.00n
.ENDS NOR3UHDV4
.SUBCKT NOR4UHDV0P7 A1 A2 A3 A4 ZN VDD VSS VNW VPW
MM3 ZN A1 VSS VPW n18 W=465.00n L=180.00n
MM5 ZN A4 VSS VPW n18 W=465.00n L=180.00n
MM9 ZN A3 VSS VPW n18 W=465.00n L=180.00n
MM1 ZN A2 VSS VPW n18 W=465.00n L=180.00n
MM2 ZN A1 net37 VNW p18 W=790.0n L=180.00n
MM0 net37 A2 net25 VNW p18 W=790.0n L=180.00n
MM4 net33 A4 VDD VNW p18 W=790.0n L=180.00n
MM8 net25 A3 net33 VNW p18 W=790.0n L=180.00n
.ENDS NOR4UHDV0P7
.SUBCKT NOR4UHDV1 A1 A2 A3 A4 ZN VDD VSS VNW VPW
MM2 ZN A1 net9 VNW p18 W=1.01u L=180.00n
MM8 net21 A3 net13 VNW p18 W=1.01u L=180.00n
MM4 net13 A4 VDD VNW p18 W=1.01u L=180.00n
MM0 net9 A2 net21 VNW p18 W=1.01u L=180.00n
MM1 ZN A2 VSS VPW n18 W=720.00n L=180.00n
MM9 ZN A3 VSS VPW n18 W=720.00n L=180.00n
MM5 ZN A4 VSS VPW n18 W=720.00n L=180.00n
MM3 ZN A1 VSS VPW n18 W=720.00n L=180.00n
.ENDS NOR4UHDV1
.SUBCKT NOR4UHDV2 A1 A2 A3 A4 ZN VDD VSS VNW VPW
MM2 ZN A1 net9 VNW p18 W=1.985u L=180.00n
MM8 net21 A3 net13 VNW p18 W=2.02u L=180.00n
MM4 net13 A4 VDD VNW p18 W=1.985u L=180.00n
MM0 net9 A2 net21 VNW p18 W=2.02u L=180.00n
MM1 ZN A2 VSS VPW n18 W=1.44u L=180.00n
MM9 ZN A3 VSS VPW n18 W=1.44u L=180.00n
MM5 ZN A4 VSS VPW n18 W=1.44u L=180.00n
MM3 ZN A1 VSS VPW n18 W=1.44u L=180.00n
.ENDS NOR4UHDV2
.SUBCKT NOR4UHDV3 A1 A2 A3 A4 ZN VDD VSS VNW VPW
MM2 ZN A1 net9 VNW p18 W=2.99u L=180.00n
MM8 net21 A3 net13 VNW p18 W=3.03u L=180.00n
MM4 net13 A4 VDD VNW p18 W=2.99u L=180.00n
MM0 net9 A2 net21 VNW p18 W=3.03u L=180.00n
MM1 ZN A2 VSS VPW n18 W=2.16u L=180.00n
MM9 ZN A3 VSS VPW n18 W=2.16u L=180.00n
MM5 ZN A4 VSS VPW n18 W=2.16u L=180.00n
MM3 ZN A1 VSS VPW n18 W=2.16u L=180.00n
.ENDS NOR4UHDV3
.SUBCKT NOR4XXBBUHDV0P7 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM10 net30 A1 net10 VPW n18 W=430.00n L=180.00n
MM3 net10 A2 VSS VPW n18 W=430.00n L=180.00n
MM1 ZN net30 VSS VPW n18 W=560.00n L=180.00n
MM5 ZN B2 VSS VPW n18 W=560.00n L=180.00n
MM9 ZN B1 VSS VPW n18 W=560.00n L=180.00n
MM11 net30 A2 VDD VNW p18 W=500.0n L=180.00n
MM2 net30 A1 VDD VNW p18 W=500.0n L=180.00n
MM8 net45 B1 net37 VNW p18 W=790.00n L=180.00n
MM4 net37 net30 VDD VNW p18 W=790.00n L=180.00n
MM0 ZN B2 net45 VNW p18 W=790.00n L=180.00n
.ENDS NOR4XXBBUHDV0P7
.SUBCKT NOR4XXBBUHDV1 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM0 ZN B2 net9 VNW p18 W=1.01u L=180.00n
MM4 net17 net18 VDD VNW p18 W=1.01u L=180.00n
MM8 net9 B1 net17 VNW p18 W=1.01u L=180.00n
MM2 net18 A1 VDD VNW p18 W=580.0n L=180.00n
MM11 net18 A2 VDD VNW p18 W=580.0n L=180.00n
MM9 ZN B1 VSS VPW n18 W=720.00n L=180.00n
MM5 ZN B2 VSS VPW n18 W=720.00n L=180.00n
MM1 ZN net18 VSS VPW n18 W=720.00n L=180.00n
MM3 net38 A2 VSS VPW n18 W=430.00n L=180.00n
MM10 net18 A1 net38 VPW n18 W=430.00n L=180.00n
.ENDS NOR4XXBBUHDV1
.SUBCKT NOR4XXBBUHDV2 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM0 ZN B2 net17 VNW p18 W=1.985u L=180.00n
MM4 net25 net10 VDD VNW p18 W=2.02u L=180.00n
MM8 net17 B1 net25 VNW p18 W=2.02u L=180.00n
MM2 net10 A1 VDD VNW p18 W=950.0n L=180.00n
MM11 net10 A2 VDD VNW p18 W=950.0n L=180.00n
MM9 ZN B1 VSS VPW n18 W=1.44u L=180.00n
MM5 ZN B2 VSS VPW n18 W=1.44u L=180.00n
MM1 ZN net10 VSS VPW n18 W=1.44u L=180.00n
MM3 net30 A2 VSS VPW n18 W=630.00n L=180.00n
MM10 net10 A1 net30 VPW n18 W=630.00n L=180.00n
.ENDS NOR4XXBBUHDV2
.SUBCKT NOR4XXBBUHDV3 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM0 ZN B2 net9 VNW p18 W=3.03u L=180.00n
MM4 net17 net18 VDD VNW p18 W=3.03u L=180.00n
MM8 net9 B1 net17 VNW p18 W=3.03u L=180.00n
MM2 net18 A1 VDD VNW p18 W=1.01u L=180.00n
MM11 net18 A2 VDD VNW p18 W=1.01u L=180.00n
MM9 ZN B1 VSS VPW n18 W=2.16u L=180.00n
MM5 ZN B2 VSS VPW n18 W=2.16u L=180.00n
MM1 ZN net18 VSS VPW n18 W=2.16u L=180.00n
MM3 net38 A2 VSS VPW n18 W=720.00n L=180.00n
MM10 net18 A1 net38 VPW n18 W=720.00n L=180.00n
.ENDS NOR4XXBBUHDV3
.SUBCKT NOR4XXBBUHDV4 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM0 ZN B2 net9 VNW p18 W=4.04u L=180.00n
MM4 net17 net18 VDD VNW p18 W=4.04u L=180.00n
MM8 net9 B1 net17 VNW p18 W=4.04u L=180.00n
MM2 net18 A1 VDD VNW p18 W=1.5u L=180.00n
MM11 net18 A2 VDD VNW p18 W=1.5u L=180.00n
MM9 ZN B1 VSS VPW n18 W=2.88u L=180.00n
MM5 ZN B2 VSS VPW n18 W=2.88u L=180.00n
MM1 ZN net18 VSS VPW n18 W=2.88u L=180.00n
MM3 net38 A2 VSS VPW n18 W=1060.00n L=180.00n
MM10 net18 A1 net38 VPW n18 W=1060.00n L=180.00n
.ENDS NOR4XXBBUHDV4
.SUBCKT OA112UHDV0P4 A1 A2 B C Z VDD VSS VNW VPW
MM8 Z net032 VSS VPW n18 W=0.28u L=180.00n
MM6 net6 C VSS VPW n18 W=0.28u L=180.00n
MM5 net21 B net6 VPW n18 W=0.28u L=180.00n
MM4 net032 A1 net21 VPW n18 W=0.28u L=180.00n
MM3 net032 A2 net21 VPW n18 W=0.28u L=180.00n
MM9 Z net032 VDD VNW p18 W=490.0n L=180.00n
MM2 net032 C VDD VNW p18 W=490.0n L=180.00n
MM1 net032 B VDD VNW p18 W=490.0n L=180.00n
MM0 net032 A1 net33 VNW p18 W=490.0n L=180.00n
MM7 net33 A2 VDD VNW p18 W=490.0n L=180.00n
.ENDS OA112UHDV0P4
.SUBCKT OA112UHDV0P7 A1 A2 B C Z VDD VSS VNW VPW
MM7 net13 A2 VDD VNW p18 W=500.0n L=180.00n
MM0 net26 A1 net13 VNW p18 W=500.0n L=180.00n
MM1 net26 B VDD VNW p18 W=500.0n L=180.00n
MM2 net26 C VDD VNW p18 W=500.0n L=180.00n
MM9 Z net26 VDD VNW p18 W=790.0n L=180.00n
MM3 net26 A2 net29 VPW n18 W=0.38u L=180.00n
MM4 net26 A1 net29 VPW n18 W=0.38u L=180.00n
MM5 net29 B net38 VPW n18 W=400.00n L=180.00n
MM6 net38 C VSS VPW n18 W=400.00n L=180.00n
MM8 Z net26 VSS VPW n18 W=560.00n L=180.00n
.ENDS OA112UHDV0P7
.SUBCKT OA112UHDV1 A1 A2 B C Z VDD VSS VNW VPW
MM7 net13 A2 VDD VNW p18 W=580.0n L=180.00n
MM0 net26 A1 net13 VNW p18 W=580.0n L=180.00n
MM1 net26 B VDD VNW p18 W=580.0n L=180.00n
MM2 net26 C VDD VNW p18 W=580.0n L=180.00n
MM9 Z net26 VDD VNW p18 W=1.01u L=180.00n
MM3 net26 A2 net29 VPW n18 W=0.38u L=180.00n
MM4 net26 A1 net29 VPW n18 W=0.38u L=180.00n
MM5 net29 B net38 VPW n18 W=400.00n L=180.00n
MM6 net38 C VSS VPW n18 W=400.00n L=180.00n
MM8 Z net26 VSS VPW n18 W=720.00n L=180.00n
.ENDS OA112UHDV1
.SUBCKT OA112UHDV2 A1 A2 B C Z VDD VSS VNW VPW
MM7 net13 A2 VDD VNW p18 W=0.92u L=180.00n
MM0 net26 A1 net13 VNW p18 W=0.92u L=180.00n
MM1 net26 B VDD VNW p18 W=0.92u L=180.00n
MM2 net26 C VDD VNW p18 W=950.0n L=180.00n
MM9 Z net26 VDD VNW p18 W=2.02u L=180.00n
MM3 net26 A2 net29 VPW n18 W=630.00n L=180.00n
MM4 net26 A1 net29 VPW n18 W=630.00n L=180.00n
MM5 net29 B net38 VPW n18 W=630.00n L=180.00n
MM6 net38 C VSS VPW n18 W=630.00n L=180.00n
MM8 Z net26 VSS VPW n18 W=1.44u L=180.00n
.ENDS OA112UHDV2
.SUBCKT OA112UHDV3 A1 A2 B C Z VDD VSS VNW VPW
MM7 net13 A2 VDD VNW p18 W=0.92u L=180.00n
MM0 net26 A1 net13 VNW p18 W=0.92u L=180.00n
MM1 net26 B VDD VNW p18 W=0.92u L=180.00n
MM2 net26 C VDD VNW p18 W=1.01u L=180.00n
MM9 Z net26 VDD VNW p18 W=3.03u L=180.00n
MM3 net26 A2 net29 VPW n18 W=720.00n L=180.00n
MM4 net26 A1 net29 VPW n18 W=720.00n L=180.00n
MM5 net29 B net38 VPW n18 W=720.00n L=180.00n
MM6 net38 C VSS VPW n18 W=720.00n L=180.00n
MM8 Z net26 VSS VPW n18 W=2.16u L=180.00n
.ENDS OA112UHDV3
.SUBCKT OA12UHDV0P4 A1 A2 B Z VDD VSS VNW VPW
MM8 Z net9 VSS VPW n18 W=0.29u L=180.00n
MM11 net12 B VSS VPW n18 W=0.26u L=180.00n
MM12 net9 A2 net12 VPW n18 W=0.28u L=180.00n
MM13 net9 A1 net12 VPW n18 W=0.26u L=180.00n
MM9 Z net9 VDD VNW p18 W=490.0n L=180.00n
MM2 net36 A2 VDD VNW p18 W=490.0n L=180.00n
MM1 net9 B VDD VNW p18 W=490.0n L=180.00n
MM10 net9 A1 net36 VNW p18 W=490.0n L=180.00n
.ENDS OA12UHDV0P4
.SUBCKT OA12UHDV0P7 A1 A2 B Z VDD VSS VNW VPW
MM10 net29 A1 net8 VNW p18 W=500.0n L=180.00n
MM1 net29 B VDD VNW p18 W=500.0n L=180.00n
MM2 net8 A2 VDD VNW p18 W=500.0n L=180.00n
MM9 Z net29 VDD VNW p18 W=790.0n L=180.00n
MM8 Z net29 VSS VPW n18 W=560.00n L=180.00n
MM13 net29 A1 net32 VPW n18 W=0.42u L=180.00n
MM12 net29 A2 net32 VPW n18 W=0.42u L=180.00n
MM11 net32 B VSS VPW n18 W=0.42u L=180.00n
.ENDS OA12UHDV0P7
.SUBCKT OA12UHDV1 A1 A2 B Z VDD VSS VNW VPW
MM10 net29 A1 net8 VNW p18 W=580.0n L=180.00n
MM1 net29 B VDD VNW p18 W=580.0n L=180.00n
MM2 net8 A2 VDD VNW p18 W=580.0n L=180.00n
MM9 Z net29 VDD VNW p18 W=1.01u L=180.00n
MM8 Z net29 VSS VPW n18 W=720.00n L=180.00n
MM13 net29 A1 net32 VPW n18 W=0.42u L=180.00n
MM12 net29 A2 net32 VPW n18 W=0.42u L=180.00n
MM11 net32 B VSS VPW n18 W=0.42u L=180.00n
.ENDS OA12UHDV1
.SUBCKT OA12UHDV2 A1 A2 B Z VDD VSS VNW VPW
MM10 net29 A1 net8 VNW p18 W=0.92u L=180.00n
MM1 net29 B VDD VNW p18 W=0.92u L=180.00n
MM2 net8 A2 VDD VNW p18 W=0.92u L=180.00n
MM9 Z net29 VDD VNW p18 W=2.02u L=180.00n
MM8 Z net29 VSS VPW n18 W=1.44u L=180.00n
MM13 net29 A1 net32 VPW n18 W=630.00n L=180.00n
MM12 net29 A2 net32 VPW n18 W=630.00n L=180.00n
MM11 net32 B VSS VPW n18 W=630.00n L=180.00n
.ENDS OA12UHDV2
.SUBCKT OA12UHDV3 A1 A2 B Z VDD VSS VNW VPW
MM10 net29 A1 net8 VNW p18 W=0.92u L=180.00n
MM1 net29 B VDD VNW p18 W=0.92u L=180.00n
MM2 net8 A2 VDD VNW p18 W=0.92u L=180.00n
MM9 Z net29 VDD VNW p18 W=3.03u L=180.00n
MM8 Z net29 VSS VPW n18 W=2.16u L=180.00n
MM13 net29 A1 net32 VPW n18 W=720.00n L=180.00n
MM12 net29 A2 net32 VPW n18 W=720.00n L=180.00n
MM11 net32 B VSS VPW n18 W=720.00n L=180.00n
.ENDS OA12UHDV3
.SUBCKT OA12UHDV4 A1 A2 B Z VDD VSS VNW VPW
MM0 Z net25 VSS VPW n18 W=2.88u L=180.00n
MM3 net25 A1 net28 VPW n18 W=1.26u L=180.00n
MM4 net25 A2 net28 VPW n18 W=1.26u L=180.00n
MM5 net28 B VSS VPW n18 W=1.26u L=180.00n
MM6 net25 A1 net52 VNW p18 W=1.84u L=180.00n
MM7 net25 B VDD VNW p18 W=1.84u L=180.00n
MM14 net52 A2 VDD VNW p18 W=1.84u L=180.00n
MM15 Z net25 VDD VNW p18 W=4.04u L=180.00n
.ENDS OA12UHDV4
.SUBCKT OA21BUHDV0P4 A1 A2 B Z VDD VSS VNW VPW
MM2 Z net17 VSS VPW n18 W=0.42u L=180.00n
MM0 Z B VSS VPW n18 W=0.42u L=180.00n
MM8 net17 A2 VSS VPW n18 W=0.42u L=180.00n
MM6 net17 A1 VSS VPW n18 W=0.42u L=180.00n
MM5 net28 net17 VDD VNW p18 W=0.5u L=180.00n
MM3 Z B net28 VNW p18 W=0.5u L=180.00n
MM1 net17 A1 net32 VNW p18 W=0.5u L=180.00n
MM4 net32 A2 VDD VNW p18 W=0.5u L=180.00n
.ENDS OA21BUHDV0P4
.SUBCKT OA21BUHDV0P7 A1 A2 B Z VDD VSS VNW VPW
MM4 net12 A2 VDD VNW p18 W=0.52u L=180.00n
MM1 net25 A1 net12 VNW p18 W=0.52u L=180.00n
MM3 Z B net16 VNW p18 W=0.81u L=180.00n
MM5 net16 net25 VDD VNW p18 W=0.81u L=180.00n
MM6 net25 A1 VSS VPW n18 W=0.48u L=180.00n
MM8 net25 A2 VSS VPW n18 W=0.48u L=180.00n
MM0 Z B VSS VPW n18 W=0.61u L=180.00n
MM2 Z net25 VSS VPW n18 W=0.61u L=180.00n
.ENDS OA21BUHDV0P7
.SUBCKT OA21BUHDV1 A1 A2 B Z VDD VSS VNW VPW
MM4 net12 A2 VDD VNW p18 W=580.0n L=180.00n
MM1 net21 A1 net12 VNW p18 W=580.0n L=180.00n
MM3 Z B net16 VNW p18 W=1.01u L=180.00n
MM5 net16 net21 VDD VNW p18 W=1.01u L=180.00n
MM8 net21 A2 VSS VPW n18 W=430.00n L=180.00n
MM6 net21 A1 VSS VPW n18 W=430.00n L=180.00n
MM0 Z B VSS VPW n18 W=720.00n L=180.00n
MM2 Z net21 VSS VPW n18 W=720.00n L=180.00n
.ENDS OA21BUHDV1
.SUBCKT OA21BUHDV2 A1 A2 B Z VDD VSS VNW VPW
MM4 net12 A2 VDD VNW p18 W=0.58u L=180.00n
MM1 net21 A1 net12 VNW p18 W=0.58u L=180.00n
MM3 Z B net16 VNW p18 W=2.02u L=180.00n
MM5 net16 net21 VDD VNW p18 W=2.02u L=180.00n
MM8 net21 A2 VSS VPW n18 W=0.43u L=180.00n
MM6 net21 A1 VSS VPW n18 W=0.43u L=180.00n
MM0 Z B VSS VPW n18 W=1.44u L=180.00n
MM2 Z net21 VSS VPW n18 W=1.44u L=180.00n
.ENDS OA21BUHDV2
.SUBCKT OA21BUHDV3 A1 A2 B Z VDD VSS VNW VPW
MM4 net12 A2 VDD VNW p18 W=1.01u L=180.00n
MM1 net21 A1 net12 VNW p18 W=1.01u L=180.00n
MM3 Z B net16 VNW p18 W=3.03u L=180.00n
MM5 net16 net21 VDD VNW p18 W=3.03u L=180.00n
MM8 net21 A2 VSS VPW n18 W=720.00n L=180.00n
MM6 net21 A1 VSS VPW n18 W=720.00n L=180.00n
MM0 Z B VSS VPW n18 W=2.16u L=180.00n
MM2 Z net21 VSS VPW n18 W=2.16u L=180.00n
.ENDS OA21BUHDV3
.SUBCKT OA221UHDV0P4 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM13 net43 B1 net31 VPW n18 W=280.00n L=180.00n
MM12 net43 B2 net31 VPW n18 W=280.00n L=180.00n
MM11 net15 C net43 VPW n18 W=280.00n L=180.00n
MM3 net31 A1 VSS VPW n18 W=280.00n L=180.00n
MM4 net31 A2 VSS VPW n18 W=280.00n L=180.00n
MM8 Z net15 VSS VPW n18 W=280.00n L=180.00n
MM10 net15 B1 net10 VNW p18 W=490.0n L=180.00n
MM7 net18 A2 VDD VNW p18 W=490.0n L=180.00n
MM0 net15 A1 net18 VNW p18 W=490.0n L=180.00n
MM1 net15 C VDD VNW p18 W=490.0n L=180.00n
MM2 net10 B2 VDD VNW p18 W=490.0n L=180.00n
MM9 Z net15 VDD VNW p18 W=490.0n L=180.00n
.ENDS OA221UHDV0P4
.SUBCKT OA221UHDV0P7 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM10 net15 B1 net10 VNW p18 W=500.0n L=180.00n
MM7 net18 A2 VDD VNW p18 W=500.0n L=180.00n
MM0 net15 A1 net18 VNW p18 W=500.0n L=180.00n
MM1 net15 C VDD VNW p18 W=500.0n L=180.00n
MM2 net10 B2 VDD VNW p18 W=500.0n L=180.00n
MM9 Z net15 VDD VNW p18 W=790.0n L=180.00n
MM13 net43 B1 net31 VPW n18 W=400.00n L=180.00n
MM12 net43 B2 net31 VPW n18 W=400.00n L=180.00n
MM11 net15 C net43 VPW n18 W=0.42u L=180.00n
MM3 net31 A1 VSS VPW n18 W=430.00n L=180.00n
MM4 net31 A2 VSS VPW n18 W=430.00n L=180.00n
MM8 Z net15 VSS VPW n18 W=560.00n L=180.00n
.ENDS OA221UHDV0P7
.SUBCKT OA221UHDV1 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM13 net23 B1 net15 VPW n18 W=0.42u L=180.00n
MM12 net23 B2 net15 VPW n18 W=0.42u L=180.00n
MM11 net43 C net23 VPW n18 W=0.42u L=180.00n
MM3 net15 A1 VSS VPW n18 W=430.00n L=180.00n
MM4 net15 A2 VSS VPW n18 W=430.00n L=180.00n
MM8 Z net43 VSS VPW n18 W=720.00n L=180.00n
MM10 net43 B1 net54 VNW p18 W=580.0n L=180.00n
MM7 net46 A2 VDD VNW p18 W=580.0n L=180.00n
MM0 net43 A1 net46 VNW p18 W=580.0n L=180.00n
MM1 net43 C VDD VNW p18 W=580.0n L=180.00n
MM2 net54 B2 VDD VNW p18 W=580.0n L=180.00n
MM9 Z net43 VDD VNW p18 W=1.01u L=180.00n
.ENDS OA221UHDV1
.SUBCKT OA221UHDV2 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM13 net23 B1 net15 VPW n18 W=630.00n L=180.00n
MM12 net23 B2 net15 VPW n18 W=630.00n L=180.00n
MM11 net43 C net23 VPW n18 W=630.00n L=180.00n
MM3 net15 A1 VSS VPW n18 W=630.00n L=180.00n
MM4 net15 A2 VSS VPW n18 W=630.00n L=180.00n
MM8 Z net43 VSS VPW n18 W=1.44u L=180.00n
MM10 net43 B1 net54 VNW p18 W=920.0n L=180.00n
MM7 net46 A2 VDD VNW p18 W=920.0n L=180.00n
MM0 net43 A1 net46 VNW p18 W=920.0n L=180.00n
MM1 net43 C VDD VNW p18 W=920.0n L=180.00n
MM2 net54 B2 VDD VNW p18 W=920.0n L=180.00n
MM9 Z net43 VDD VNW p18 W=2.02u L=180.00n
.ENDS OA221UHDV2
.SUBCKT OA221UHDV3 A1 A2 B1 B2 C Z VDD VSS VNW VPW
MM10 net101 B1 net112 VNW p18 W=1.54u L=180.00n
MM7 net104 A2 VDD VNW p18 W=1.74u L=180.00n
MM0 net101 A1 net104 VNW p18 W=1.74u L=180.00n
MM1 net101 C VDD VNW p18 W=1.74u L=180.00n
MM2 net112 B2 VDD VNW p18 W=1.54u L=180.00n
MM9 Z net101 VDD VNW p18 W=3.03u L=180.00n
MM13 net129 B1 net121 VPW n18 W=1.12u L=180.00n
MM12 net129 B2 net121 VPW n18 W=1.12u L=180.00n
MM11 net101 C net129 VPW n18 W=1.26u L=180.00n
MM3 net121 A1 VSS VPW n18 W=1.26u L=180.00n
MM4 net121 A2 VSS VPW n18 W=1.26u L=180.00n
MM8 Z net101 VSS VPW n18 W=2.16u L=180.00n
.ENDS OA221UHDV3
.SUBCKT OA222UHDV0P4 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM8 Z net40 VSS VPW n18 W=280.00n L=180.00n
MM4 net48 C1 VSS VPW n18 W=280.00n L=180.00n
MM3 net48 C2 VSS VPW n18 W=280.00n L=180.00n
MM6 net40 A2 net52 VPW n18 W=280.00n L=180.00n
MM12 net52 B2 net48 VPW n18 W=280.00n L=180.00n
MM13 net52 B1 net48 VPW n18 W=280.00n L=180.00n
MM11 net40 A1 net52 VPW n18 W=280.00n L=180.00n
MM5 net40 A2 net11 VNW p18 W=490.0n L=180.00n
MM9 Z net40 VDD VNW p18 W=490.0n L=180.00n
MM2 net35 B2 VDD VNW p18 W=490.0n L=180.00n
MM1 net11 A1 VDD VNW p18 W=490.0n L=180.00n
MM0 net40 C2 net27 VNW p18 W=490.0n L=180.00n
MM7 net27 C1 VDD VNW p18 W=490.0n L=180.00n
MM10 net40 B1 net35 VNW p18 W=490.0n L=180.00n
.ENDS OA222UHDV0P4
.SUBCKT OA222UHDV0P7 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM8 Z net40 VSS VPW n18 W=560.00n L=180.00n
MM4 net48 C1 VSS VPW n18 W=400.00n L=180.00n
MM3 net48 C2 VSS VPW n18 W=400.00n L=180.00n
MM6 net40 A2 net52 VPW n18 W=400.00n L=180.00n
MM12 net52 B2 net48 VPW n18 W=400.00n L=180.00n
MM13 net52 B1 net48 VPW n18 W=400.00n L=180.00n
MM11 net40 A1 net52 VPW n18 W=400.00n L=180.00n
MM5 net40 A2 net11 VNW p18 W=500.0n L=180.00n
MM9 Z net40 VDD VNW p18 W=790.0n L=180.00n
MM2 net35 B2 VDD VNW p18 W=500.0n L=180.00n
MM1 net11 A1 VDD VNW p18 W=500.0n L=180.00n
MM0 net40 C2 net27 VNW p18 W=500.0n L=180.00n
MM7 net27 C1 VDD VNW p18 W=500.0n L=180.00n
MM10 net40 B1 net35 VNW p18 W=500.0n L=180.00n
.ENDS OA222UHDV0P7
.SUBCKT OA222UHDV1 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM5 net40 A2 net11 VNW p18 W=580.0n L=180.00n
MM9 Z net40 VDD VNW p18 W=1.01u L=180.00n
MM2 net35 B2 VDD VNW p18 W=580.0n L=180.00n
MM1 net11 A1 VDD VNW p18 W=580.0n L=180.00n
MM0 net40 C2 net27 VNW p18 W=580.0n L=180.00n
MM7 net27 C1 VDD VNW p18 W=580.0n L=180.00n
MM10 net40 B1 net35 VNW p18 W=580.0n L=180.00n
MM8 Z net40 VSS VPW n18 W=720.00n L=180.00n
MM4 net48 C1 VSS VPW n18 W=0.42u L=180.00n
MM3 net48 C2 VSS VPW n18 W=0.42u L=180.00n
MM6 net40 A2 net52 VPW n18 W=0.38u L=180.00n
MM12 net52 B2 net48 VPW n18 W=0.38u L=180.00n
MM13 net52 B1 net48 VPW n18 W=0.38u L=180.00n
MM11 net40 A1 net52 VPW n18 W=0.38u L=180.00n
.ENDS OA222UHDV1
.SUBCKT OA222UHDV2 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM8 Z net40 VSS VPW n18 W=1.44u L=180.00n
MM4 net48 C1 VSS VPW n18 W=660.00n L=180.00n
MM3 net48 C2 VSS VPW n18 W=660.00n L=180.00n
MM6 net40 A2 net52 VPW n18 W=620.00n L=180.00n
MM12 net52 B2 net48 VPW n18 W=620.00n L=180.00n
MM13 net52 B1 net48 VPW n18 W=620.00n L=180.00n
MM11 net40 A1 net52 VPW n18 W=620.00n L=180.00n
MM5 net40 A2 net11 VNW p18 W=950.00n L=180.00n
MM9 Z net40 VDD VNW p18 W=2.02u L=180.00n
MM2 net35 B2 VDD VNW p18 W=950.00n L=180.00n
MM1 net11 A1 VDD VNW p18 W=950.00n L=180.00n
MM0 net40 C2 net27 VNW p18 W=1.01u L=180.00n
MM7 net27 C1 VDD VNW p18 W=1.01u L=180.00n
MM10 net40 B1 net35 VNW p18 W=950.00n L=180.00n
.ENDS OA222UHDV2
.SUBCKT OA222UHDV3 A1 A2 B1 B2 C1 C2 Z VDD VSS VNW VPW
MM8 Z net40 VSS VPW n18 W=2.16u L=180.00n
MM4 net48 C1 VSS VPW n18 W=1.14u L=180.00n
MM3 net48 C2 VSS VPW n18 W=1u L=180.00n
MM6 net40 A2 net52 VPW n18 W=1.14u L=180.00n
MM12 net52 B2 net48 VPW n18 W=1.14u L=180.00n
MM13 net52 B1 net48 VPW n18 W=1u L=180.00n
MM11 net40 A1 net52 VPW n18 W=1.14u L=180.00n
MM5 net40 A2 net11 VNW p18 W=1.74u L=180.00n
MM9 Z net40 VDD VNW p18 W=3.03u L=180.00n
MM2 net35 B2 VDD VNW p18 W=1.74u L=180.00n
MM1 net11 A1 VDD VNW p18 W=1.74u L=180.00n
MM0 net40 C2 net27 VNW p18 W=1.54u L=180.00n
MM7 net27 C1 VDD VNW p18 W=1.74u L=180.00n
MM10 net40 B1 net35 VNW p18 W=1.54u L=180.00n
.ENDS OA222UHDV3
.SUBCKT OA22UHDV0P4 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM8 Z net18 VSS VPW n18 W=280.00n L=180.00n
MM13 net14 B1 VSS VPW n18 W=280.00n L=180.00n
MM12 net14 B2 VSS VPW n18 W=280.00n L=180.00n
MM6 net18 A1 net14 VPW n18 W=280.00n L=180.00n
MM11 net18 A2 net14 VPW n18 W=280.00n L=180.00n
MM10 net18 B1 net37 VNW p18 W=490.0n L=180.00n
MM1 net33 A2 VDD VNW p18 W=490.0n L=180.00n
MM2 net37 B2 VDD VNW p18 W=490.0n L=180.00n
MM9 Z net18 VDD VNW p18 W=490.0n L=180.00n
MM5 net18 A1 net33 VNW p18 W=490.0n L=180.00n
.ENDS OA22UHDV0P4
.SUBCKT OA22UHDV0P7 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM8 Z net18 VSS VPW n18 W=560.00n L=180.00n
MM13 net14 B1 VSS VPW n18 W=430.00n L=180.00n
MM12 net14 B2 VSS VPW n18 W=430.00n L=180.00n
MM6 net18 A1 net14 VPW n18 W=430.00n L=180.00n
MM11 net18 A2 net14 VPW n18 W=430.00n L=180.00n
MM10 net18 B1 net37 VNW p18 W=500.0n L=180.00n
MM1 net33 A2 VDD VNW p18 W=500.0n L=180.00n
MM2 net37 B2 VDD VNW p18 W=500.0n L=180.00n
MM9 Z net18 VDD VNW p18 W=790.0n L=180.00n
MM5 net18 A1 net33 VNW p18 W=500.0n L=180.00n
.ENDS OA22UHDV0P7
.SUBCKT OA22UHDV1 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM8 Z net18 VSS VPW n18 W=720.00n L=180.00n
MM13 net14 B1 VSS VPW n18 W=0.38u L=180.00n
MM12 net14 B2 VSS VPW n18 W=0.38u L=180.00n
MM6 net18 A1 net14 VPW n18 W=0.38u L=180.00n
MM11 net18 A2 net14 VPW n18 W=0.38u L=180.00n
MM10 net18 B1 net37 VNW p18 W=580.0n L=180.00n
MM1 net33 A2 VDD VNW p18 W=580.0n L=180.00n
MM2 net37 B2 VDD VNW p18 W=580.0n L=180.00n
MM9 Z net18 VDD VNW p18 W=1.01u L=180.00n
MM5 net18 A1 net33 VNW p18 W=580.0n L=180.00n
.ENDS OA22UHDV1
.SUBCKT OA22UHDV2 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM9 Z net30 VDD VNW p18 W=2.02u L=180.00n
MM2 net17 B2 VDD VNW p18 W=0.925u L=180.00n
MM10 net30 B1 net17 VNW p18 W=0.925u L=180.00n
MM5 net30 A1 net21 VNW p18 W=0.925u L=180.00n
MM1 net21 A2 VDD VNW p18 W=0.925u L=180.00n
MM8 Z net30 VSS VPW n18 W=1.44u L=180.00n
MM6 net30 A1 net33 VPW n18 W=0.63u L=180.00n
MM12 net33 B2 VSS VPW n18 W=630.00n L=180.00n
MM11 net30 A2 net33 VPW n18 W=600.00n L=180.00n
MM13 net33 B1 VSS VPW n18 W=630.00n L=180.00n
.ENDS OA22UHDV2
.SUBCKT OA22UHDV3 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM8 Z net18 VSS VPW n18 W=2.16u L=180.00n
MM13 net14 B1 VSS VPW n18 W=1.14u L=180.00n
MM12 net14 B2 VSS VPW n18 W=1.14u L=180.00n
MM6 net18 A1 net14 VPW n18 W=1.14u L=180.00n
MM11 net18 A2 net14 VPW n18 W=1.14u L=180.00n
MM10 net18 B1 net37 VNW p18 W=1.74u L=180.00n
MM1 net33 A2 VDD VNW p18 W=1.74u L=180.00n
MM2 net37 B2 VDD VNW p18 W=1.74u L=180.00n
MM9 Z net18 VDD VNW p18 W=3.03u L=180.00n
MM5 net18 A1 net33 VNW p18 W=1.74u L=180.00n
.ENDS OA22UHDV3
.SUBCKT OA22UHDV4 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM8 Z net18 VSS VPW n18 W=2.88u L=180.00n
MM13 net14 B1 VSS VPW n18 W=1.28u L=180.00n
MM12 net14 B2 VSS VPW n18 W=1.28u L=180.00n
MM6 net18 A1 net14 VPW n18 W=1.2u L=180.00n
MM11 net18 A2 net14 VPW n18 W=1.2u L=180.00n
MM10 net18 B1 net37 VNW p18 W=1.95u L=180.00n
MM1 net33 A2 VDD VNW p18 W=1.86u L=180.00n
MM2 net37 B2 VDD VNW p18 W=1.95u L=180.00n
MM9 Z net18 VDD VNW p18 W=4.04u L=180.00n
MM5 net18 A1 net33 VNW p18 W=1.86u L=180.00n
.ENDS OA22UHDV4
.SUBCKT OA22UHDV6 A1 A2 B1 B2 Z VDD VSS VNW VPW
MM8 Z net18 VSS VPW n18 W=4.42u L=180.00n
MM13 net14 B1 VSS VPW n18 W=2.28u L=180.00n
MM12 net14 B2 VSS VPW n18 W=2.28u L=180.00n
MM6 net18 A1 net14 VPW n18 W=2.28u L=180.00n
MM11 net18 A2 net14 VPW n18 W=2.28u L=180.00n
MM10 net18 B1 net37 VNW p18 W=3.48u L=180.00n
MM1 net33 A2 VDD VNW p18 W=3.48u L=180.00n
MM2 net37 B2 VDD VNW p18 W=3.48u L=180.00n
MM9 Z net18 VDD VNW p18 W=6.06u L=180.00n
MM5 net18 A1 net33 VNW p18 W=3.48u L=180.00n
.ENDS OA22UHDV6
.SUBCKT OA31UHDV0P4 A1 A2 A3 B Z VDD VSS VNW VPW
MM0 net21 A3 VDD VNW p18 W=490.0n L=180.00n
MM10 net6 A1 net17 VNW p18 W=490.0n L=180.00n
MM1 net6 B VDD VNW p18 W=490.0n L=180.00n
MM2 net17 A2 net21 VNW p18 W=490.0n L=180.00n
MM9 Z net6 VDD VNW p18 W=490.0n L=180.00n
MM3 net30 A2 VSS VPW n18 W=0.28u L=180.00n
MM8 Z net6 VSS VPW n18 W=0.28u L=180.00n
MM13 net30 A1 VSS VPW n18 W=0.28u L=180.00n
MM12 net30 A3 VSS VPW n18 W=0.28u L=180.00n
MM11 net6 B net30 VPW n18 W=0.28u L=180.00n
.ENDS OA31UHDV0P4
.SUBCKT OA31UHDV0P7 A1 A2 A3 B Z VDD VSS VNW VPW
MM8 Z net42 VSS VPW n18 W=500.00n L=180.00n
MM11 net42 B net18 VPW n18 W=300.00n L=180.00n
MM13 net18 A1 VSS VPW n18 W=300.00n L=180.00n
MM12 net18 A3 VSS VPW n18 W=300.00n L=180.00n
MM3 net18 A2 VSS VPW n18 W=300.00n L=180.00n
MM9 Z net42 VDD VNW p18 W=700.0n L=180.00n
MM2 net37 A2 net33 VNW p18 W=400.0n L=180.00n
MM10 net42 A1 net37 VNW p18 W=400.0n L=180.00n
MM0 net33 A3 VDD VNW p18 W=400.0n L=180.00n
MM1 net42 B VDD VNW p18 W=400.0n L=180.00n
.ENDS OA31UHDV0P7
.SUBCKT OA31UHDV1 A1 A2 A3 B Z VDD VSS VNW VPW
MM8 Z net42 VSS VPW n18 W=720.00n L=180.00n
MM11 net42 B net18 VPW n18 W=0.44u L=180.00n
MM13 net18 A1 VSS VPW n18 W=0.44u L=180.00n
MM12 net18 A3 VSS VPW n18 W=0.44u L=180.00n
MM3 net18 A2 VSS VPW n18 W=0.44u L=180.00n
MM9 Z net42 VDD VNW p18 W=1.01u L=180.00n
MM2 net37 A2 net33 VNW p18 W=580.0n L=180.00n
MM10 net42 A1 net37 VNW p18 W=580.0n L=180.00n
MM0 net33 A3 VDD VNW p18 W=580.0n L=180.00n
MM1 net42 B VDD VNW p18 W=580.0n L=180.00n
.ENDS OA31UHDV1
.SUBCKT OA31UHDV2 A1 A2 A3 B Z VDD VSS VNW VPW
MM8 Z net42 VSS VPW n18 W=1.44u L=180.00n
MM11 net42 B net18 VPW n18 W=720.00n L=180.00n
MM13 net18 A1 VSS VPW n18 W=720.00n L=180.00n
MM12 net18 A3 VSS VPW n18 W=720.00n L=180.00n
MM3 net18 A2 VSS VPW n18 W=720.00n L=180.00n
MM9 Z net42 VDD VNW p18 W=2.02u L=180.00n
MM2 net37 A2 net33 VNW p18 W=950.00n L=180.00n
MM10 net42 A1 net37 VNW p18 W=950.00n L=180.00n
MM0 net33 A3 VDD VNW p18 W=950.00n L=180.00n
MM1 net42 B VDD VNW p18 W=950.00n L=180.00n
.ENDS OA31UHDV2
.SUBCKT OA32UHDV0P7 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM0 net26 A3 VDD VNW p18 W=500.0n L=180.00n
MM5 net43 A1 net18 VNW p18 W=500.0n L=180.00n
MM9 Z net43 VDD VNW p18 W=790.0n L=180.00n
MM2 net30 B2 VDD VNW p18 W=500.0n L=180.00n
MM1 net18 A2 net26 VNW p18 W=500.0n L=180.00n
MM10 net43 B1 net30 VNW p18 W=500.0n L=180.00n
MM11 net43 A2 net47 VPW n18 W=430.00n L=180.00n
MM6 net43 A1 net47 VPW n18 W=430.00n L=180.00n
MM12 net47 B2 VSS VPW n18 W=430.00n L=180.00n
MM13 net47 B1 VSS VPW n18 W=430.00n L=180.00n
MM8 Z net43 VSS VPW n18 W=560.00n L=180.00n
MM3 net43 A3 net47 VPW n18 W=430.00n L=180.00n
.ENDS OA32UHDV0P7
.SUBCKT OA32UHDV1 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM13 net11 B1 VSS VPW n18 W=430.00n L=180.00n
MM12 net11 B2 VSS VPW n18 W=430.00n L=180.00n
MM6 net15 A1 net11 VPW n18 W=430.00n L=180.00n
MM11 net15 A2 net11 VPW n18 W=430.00n L=180.00n
MM8 Z net15 VSS VPW n18 W=720.00n L=180.00n
MM3 net15 A3 net11 VPW n18 W=430.00n L=180.00n
MM10 net15 B1 net34 VNW p18 W=580.0n L=180.00n
MM1 net46 A2 net38 VNW p18 W=580.0n L=180.00n
MM2 net34 B2 VDD VNW p18 W=580.0n L=180.00n
MM5 net15 A1 net46 VNW p18 W=580.0n L=180.00n
MM0 net38 A3 VDD VNW p18 W=580.0n L=180.00n
MM9 Z net15 VDD VNW p18 W=1.01u L=180.00n
.ENDS OA32UHDV1
.SUBCKT OA32UHDV2 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM9 Z net43 VDD VNW p18 W=2.02u L=180.00n
MM0 net26 A3 VDD VNW p18 W=950.0n L=180.00n
MM5 net43 A1 net18 VNW p18 W=0.92u L=180.00n
MM2 net30 B2 VDD VNW p18 W=950.0n L=180.00n
MM1 net18 A2 net26 VNW p18 W=0.92u L=180.00n
MM10 net43 B1 net30 VNW p18 W=950.0n L=180.00n
MM3 net43 A3 net47 VPW n18 W=630.00n L=180.00n
MM8 Z net43 VSS VPW n18 W=1.44u L=180.00n
MM11 net43 A2 net47 VPW n18 W=630.00n L=180.00n
MM6 net43 A1 net47 VPW n18 W=630.00n L=180.00n
MM12 net47 B2 VSS VPW n18 W=630.00n L=180.00n
MM13 net47 B1 VSS VPW n18 W=630.00n L=180.00n
.ENDS OA32UHDV2
.SUBCKT OA32UHDV3 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM13 net11 B1 VSS VPW n18 W=720.00n L=180.00n
MM12 net11 B2 VSS VPW n18 W=720.00n L=180.00n
MM6 net15 A1 net11 VPW n18 W=720.00n L=180.00n
MM11 net15 A2 net11 VPW n18 W=720.00n L=180.00n
MM8 Z net15 VSS VPW n18 W=2.16u L=180.00n
MM3 net15 A3 net11 VPW n18 W=720.00n L=180.00n
MM10 net15 B1 net34 VNW p18 W=1.01u L=180.00n
MM1 net46 A2 net38 VNW p18 W=0.92u L=180.00n
MM2 net34 B2 VDD VNW p18 W=1.01u L=180.00n
MM5 net15 A1 net46 VNW p18 W=0.92u L=180.00n
MM0 net38 A3 VDD VNW p18 W=1.01u L=180.00n
MM9 Z net15 VDD VNW p18 W=3.03u L=180.00n
.ENDS OA32UHDV3
.SUBCKT OA32UHDV4 A1 A2 A3 B1 B2 Z VDD VSS VNW VPW
MM9 Z net43 VDD VNW p18 W=4.04u L=180.00n
MM0 net26 A3 VDD VNW p18 W=1.49u L=180.00n
MM5 net43 A1 net18 VNW p18 W=1.49u L=180.00n
MM2 net30 B2 VDD VNW p18 W=1.49u L=180.00n
MM1 net18 A2 net26 VNW p18 W=1.49u L=180.00n
MM10 net43 B1 net30 VNW p18 W=1.49u L=180.00n
MM3 net43 A3 net47 VPW n18 W=1060.00n L=180.00n
MM8 Z net43 VSS VPW n18 W=2.88u L=180.00n
MM11 net43 A2 net47 VPW n18 W=1060.00n L=180.00n
MM6 net43 A1 net47 VPW n18 W=1060.00n L=180.00n
MM12 net47 B2 VSS VPW n18 W=1060.00n L=180.00n
MM13 net47 B1 VSS VPW n18 W=1060.00n L=180.00n
.ENDS OA32UHDV4
.SUBCKT OA33UHDV0P7 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM7 net24 B3 VSS VPW n18 W=430.00n L=180.00n
MM3 net28 A3 net24 VPW n18 W=0.44u L=180.00n
MM8 Z net28 VSS VPW n18 W=560.00n L=180.00n
MM13 net24 B1 VSS VPW n18 W=430.00n L=180.00n
MM12 net24 B2 VSS VPW n18 W=430.00n L=180.00n
MM6 net28 A1 net24 VPW n18 W=430.00n L=180.00n
MM11 net28 A2 net24 VPW n18 W=0.44u L=180.00n
MM4 net51 B3 VDD VNW p18 W=500.0n L=180.00n
MM10 net28 B1 net43 VNW p18 W=500.0n L=180.00n
MM1 net59 A2 net47 VNW p18 W=500.0n L=180.00n
MM2 net43 B2 net51 VNW p18 W=500.0n L=180.00n
MM9 Z net28 VDD VNW p18 W=790.0n L=180.00n
MM5 net28 A1 net59 VNW p18 W=500.0n L=180.00n
MM0 net47 A3 VDD VNW p18 W=500.0n L=180.00n
.ENDS OA33UHDV0P7
.SUBCKT OA33UHDV1 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM0 net27 A3 VDD VNW p18 W=580.0n L=180.00n
MM5 net40 A1 net15 VNW p18 W=580.0n L=180.00n
MM9 Z net40 VDD VNW p18 W=1.01u L=180.00n
MM2 net31 B2 net23 VNW p18 W=580.0n L=180.00n
MM1 net15 A2 net27 VNW p18 W=580.0n L=180.00n
MM10 net40 B1 net31 VNW p18 W=580.0n L=180.00n
MM4 net23 B3 VDD VNW p18 W=580.0n L=180.00n
MM11 net40 A2 net44 VPW n18 W=430.00n L=180.00n
MM6 net40 A1 net44 VPW n18 W=430.00n L=180.00n
MM12 net44 B2 VSS VPW n18 W=430.00n L=180.00n
MM13 net44 B1 VSS VPW n18 W=430.00n L=180.00n
MM8 Z net40 VSS VPW n18 W=720.00n L=180.00n
MM3 net40 A3 net44 VPW n18 W=430.00n L=180.00n
MM7 net44 B3 VSS VPW n18 W=430.00n L=180.00n
.ENDS OA33UHDV1
.SUBCKT OA33UHDV2 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM7 net24 B3 VSS VPW n18 W=630.00n L=180.00n
MM3 net28 A3 net24 VPW n18 W=630.00n L=180.00n
MM8 Z net28 VSS VPW n18 W=1.44u L=180.00n
MM13 net24 B1 VSS VPW n18 W=630.00n L=180.00n
MM12 net24 B2 VSS VPW n18 W=630.00n L=180.00n
MM6 net28 A1 net24 VPW n18 W=630.00n L=180.00n
MM11 net28 A2 net24 VPW n18 W=630.00n L=180.00n
MM4 net51 B3 VDD VNW p18 W=950.0n L=180.00n
MM10 net28 B1 net43 VNW p18 W=0.92u L=180.00n
MM1 net59 A2 net47 VNW p18 W=0.92u L=180.00n
MM2 net43 B2 net51 VNW p18 W=950.0n L=180.00n
MM9 Z net28 VDD VNW p18 W=2.02u L=180.00n
MM5 net28 A1 net59 VNW p18 W=0.92u L=180.00n
MM0 net47 A3 VDD VNW p18 W=950.0n L=180.00n
.ENDS OA33UHDV2
.SUBCKT OA33UHDV3 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM0 net27 A3 VDD VNW p18 W=1.01u L=180.00n
MM5 net40 A1 net15 VNW p18 W=0.92u L=180.00n
MM9 Z net40 VDD VNW p18 W=3.03u L=180.00n
MM2 net31 B2 net23 VNW p18 W=1.01u L=180.00n
MM1 net15 A2 net27 VNW p18 W=0.92u L=180.00n
MM10 net40 B1 net31 VNW p18 W=0.92u L=180.00n
MM4 net23 B3 VDD VNW p18 W=1.01u L=180.00n
MM11 net40 A2 net44 VPW n18 W=720.00n L=180.00n
MM6 net40 A1 net44 VPW n18 W=720.00n L=180.00n
MM12 net44 B2 VSS VPW n18 W=720.00n L=180.00n
MM13 net44 B1 VSS VPW n18 W=720.00n L=180.00n
MM8 Z net40 VSS VPW n18 W=2.16u L=180.00n
MM3 net40 A3 net44 VPW n18 W=720.00n L=180.00n
MM7 net44 B3 VSS VPW n18 W=720.00n L=180.00n
.ENDS OA33UHDV3
.SUBCKT OA33UHDV4 A1 A2 A3 B1 B2 B3 Z VDD VSS VNW VPW
MM7 net24 B3 VSS VPW n18 W=1060.00n L=180.00n
MM3 net28 A3 net24 VPW n18 W=1060.00n L=180.00n
MM8 Z net28 VSS VPW n18 W=2.88u L=180.00n
MM13 net24 B1 VSS VPW n18 W=1060.00n L=180.00n
MM12 net24 B2 VSS VPW n18 W=1060.00n L=180.00n
MM6 net28 A1 net24 VPW n18 W=1060.00n L=180.00n
MM11 net28 A2 net24 VPW n18 W=1060.00n L=180.00n
MM4 net51 B3 VDD VNW p18 W=1.49u L=180.00n
MM10 net28 B1 net43 VNW p18 W=1.49u L=180.00n
MM1 net59 A2 net47 VNW p18 W=1.49u L=180.00n
MM2 net43 B2 net51 VNW p18 W=1.49u L=180.00n
MM9 Z net28 VDD VNW p18 W=4.04u L=180.00n
MM5 net28 A1 net59 VNW p18 W=1.49u L=180.00n
MM0 net47 A3 VDD VNW p18 W=1.49u L=180.00n
.ENDS OA33UHDV4
.SUBCKT OAI211UHDV0P4 A1 A2 B C ZN VDD VSS VNW VPW
MM7 net13 A2 VDD VNW p18 W=0.48u L=180.00n
MM0 ZN A1 net13 VNW p18 W=0.48u L=180.00n
MM1 ZN B VDD VNW p18 W=0.48u L=180.00n
MM2 ZN C VDD VNW p18 W=0.48u L=180.00n
MM3 net26 A2 VSS VPW n18 W=0.28u L=180.00n
MM4 net26 A1 VSS VPW n18 W=0.28u L=180.00n
MM5 ZN B net38 VPW n18 W=0.28u L=180.00n
MM6 net38 C net26 VPW n18 W=0.28u L=180.00n
.ENDS OAI211UHDV0P4
.SUBCKT OAI211UHDV0P7 A1 A2 B C ZN VDD VSS VNW VPW
MM6 net6 C net18 VPW n18 W=560.00n L=180.00n
MM5 ZN B net6 VPW n18 W=560.00n L=180.00n
MM4 net18 A1 VSS VPW n18 W=0.56u L=180.00n
MM3 net18 A2 VSS VPW n18 W=0.535u L=180.00n
MM2 ZN C VDD VNW p18 W=540.0n L=180.00n
MM1 ZN B VDD VNW p18 W=540.0n L=180.00n
MM0 ZN A1 net33 VNW p18 W=790.0n L=180.00n
MM7 net33 A2 VDD VNW p18 W=790.0n L=180.00n
.ENDS OAI211UHDV0P7
.SUBCKT OAI211UHDV1 A1 A2 B C ZN VDD VSS VNW VPW
MM6 net6 C net18 VPW n18 W=720.00n L=180.00n
MM5 ZN B net6 VPW n18 W=720.00n L=180.00n
MM4 net18 A1 VSS VPW n18 W=720.00n L=180.00n
MM3 net18 A2 VSS VPW n18 W=720.00n L=180.00n
MM2 ZN C VDD VNW p18 W=1.01u L=180.00n
MM1 ZN B VDD VNW p18 W=1.01u L=180.00n
MM0 ZN A1 net33 VNW p18 W=1.01u L=180.00n
MM7 net33 A2 VDD VNW p18 W=1.01u L=180.00n
.ENDS OAI211UHDV1
.SUBCKT OAI211UHDV2 A1 A2 B C ZN VDD VSS VNW VPW
MM6 net6 C net18 VPW n18 W=1.44u L=180.00n
MM5 ZN B net6 VPW n18 W=1.55u L=180.00n
MM4 net18 A1 VSS VPW n18 W=1.44u L=180.00n
MM3 net18 A2 VSS VPW n18 W=1.44u L=180.00n
MM2 ZN C VDD VNW p18 W=1.49u L=180.00n
MM1 ZN B VDD VNW p18 W=1.49u L=180.00n
MM0 ZN A1 net33 VNW p18 W=1.95u L=180.00n
MM7 net33 A2 VDD VNW p18 W=2.02u L=180.00n
.ENDS OAI211UHDV2
.SUBCKT OAI211UHDV3 A1 A2 B C ZN VDD VSS VNW VPW
MM6 net6 C net18 VPW n18 W=2.16u L=180.00n
MM5 ZN B net6 VPW n18 W=2.16u L=180.00n
MM4 net18 A1 VSS VPW n18 W=2.16u L=180.00n
MM3 net18 A2 VSS VPW n18 W=2.16u L=180.00n
MM2 ZN C VDD VNW p18 W=1.9u L=180.00n
MM1 ZN B VDD VNW p18 W=1.47u L=180.00n
MM0 ZN A1 net33 VNW p18 W=2.96u L=180.00n
MM7 net33 A2 VDD VNW p18 W=3.03u L=180.00n
.ENDS OAI211UHDV3
.SUBCKT OAI21BUHDV0P4 A B1 B2 ZN VDD VSS VNW VPW
MM10 ZN B1 net8 VNW p18 W=490.0n L=180.00n
MM1 ZN net33 VDD VNW p18 W=490.0n L=180.00n
MM2 net8 B2 VDD VNW p18 W=490.0n L=180.00n
MM3 net33 A VDD VNW p18 W=490.0n L=180.00n
MM0 ZN net33 net29 VPW n18 W=420.00n L=180.00n
MM13 net29 B1 VSS VPW n18 W=420.00n L=180.00n
MM12 net29 B2 VSS VPW n18 W=420.00n L=180.00n
MM4 net33 A VSS VPW n18 W=430.00n L=180.00n
.ENDS OAI21BUHDV0P4
.SUBCKT OAI21BUHDV0P7 A B1 B2 ZN VDD VSS VNW VPW
MM4 net5 A VSS VPW n18 W=430.00n L=180.00n
MM12 net9 B2 VSS VPW n18 W=560.00n L=180.00n
MM13 net9 B1 VSS VPW n18 W=560.00n L=180.00n
MM0 ZN net5 net9 VPW n18 W=560.00n L=180.00n
MM3 net5 A VDD VNW p18 W=500.0n L=180.00n
MM2 net36 B2 VDD VNW p18 W=790.0n L=180.00n
MM1 ZN net5 VDD VNW p18 W=790.0n L=180.00n
MM10 ZN B1 net36 VNW p18 W=790.0n L=180.00n
.ENDS OAI21BUHDV0P7
.SUBCKT OAI21BUHDV1 A B1 B2 ZN VDD VSS VNW VPW
MM10 ZN B1 net8 VNW p18 W=1.01u L=180.00n
MM1 ZN net33 VDD VNW p18 W=1.01u L=180.00n
MM2 net8 B2 VDD VNW p18 W=1.01u L=180.00n
MM3 net33 A VDD VNW p18 W=580.0n L=180.00n
MM0 ZN net33 net29 VPW n18 W=720.00n L=180.00n
MM13 net29 B1 VSS VPW n18 W=720.00n L=180.00n
MM12 net29 B2 VSS VPW n18 W=720.00n L=180.00n
MM4 net33 A VSS VPW n18 W=430.00n L=180.00n
.ENDS OAI21BUHDV1
.SUBCKT OAI21BUHDV2 A B1 B2 ZN VDD VSS VNW VPW
MM4 net5 A VSS VPW n18 W=630.00n L=180.00n
MM12 net9 B2 VSS VPW n18 W=1.415u L=180.00n
MM13 net9 B1 VSS VPW n18 W=1.39u L=180.00n
MM0 ZN net5 net9 VPW n18 W=1.44u L=180.00n
MM3 net5 A VDD VNW p18 W=950.0n L=180.00n
MM2 net36 B2 VDD VNW p18 W=1.985u L=180.00n
MM1 ZN net5 VDD VNW p18 W=1.9u L=180.00n
MM10 ZN B1 net36 VNW p18 W=2.02u L=180.00n
.ENDS OAI21BUHDV2
.SUBCKT OAI21UHDV0P4 A1 A2 B ZN VDD VSS VNW VPW
MM10 ZN A1 net8 VNW p18 W=490.0n L=180.00n
MM1 ZN B VDD VNW p18 W=490.0n L=180.00n
MM2 net8 A2 VDD VNW p18 W=490.0n L=180.00n
MM0 ZN B net17 VPW n18 W=0.28u L=180.00n
MM13 net17 A1 VSS VPW n18 W=0.28u L=180.00n
MM12 net17 A2 VSS VPW n18 W=0.28u L=180.00n
.ENDS OAI21UHDV0P4
.SUBCKT OAI21UHDV0P7 A1 A2 B ZN VDD VSS VNW VPW
MM0 ZN B net13 VPW n18 W=560.00n L=180.00n
MM13 net13 A1 VSS VPW n18 W=560.00n L=180.00n
MM12 net13 A2 VSS VPW n18 W=560.00n L=180.00n
MM2 net28 A2 VDD VNW p18 W=790.0n L=180.00n
MM1 ZN B VDD VNW p18 W=790.0n L=180.00n
MM10 ZN A1 net28 VNW p18 W=790.0n L=180.00n
.ENDS OAI21UHDV0P7
.SUBCKT OAI21UHDV1 A1 A2 B ZN VDD VSS VNW VPW
MM0 ZN B net13 VPW n18 W=720.00n L=180.00n
MM13 net13 A1 VSS VPW n18 W=720.00n L=180.00n
MM12 net13 A2 VSS VPW n18 W=720.00n L=180.00n
MM2 net28 A2 VDD VNW p18 W=1.01u L=180.00n
MM1 ZN B VDD VNW p18 W=1.01u L=180.00n
MM10 ZN A1 net28 VNW p18 W=1.01u L=180.00n
.ENDS OAI21UHDV1
.SUBCKT OAI21UHDV2 A1 A2 B ZN VDD VSS VNW VPW
MM0 ZN B net13 VPW n18 W=1.44u L=180.00n
MM13 net13 A1 VSS VPW n18 W=1.44u L=180.00n
MM12 net13 A2 VSS VPW n18 W=1.44u L=180.00n
MM2 net28 A2 VDD VNW p18 W=2.02u L=180.00n
MM1 ZN B VDD VNW p18 W=1.85u L=180.00n
MM10 ZN A1 net28 VNW p18 W=2.02u L=180.00n
.ENDS OAI21UHDV2
.SUBCKT OAI21UHDV3 A1 A2 B ZN VDD VSS VNW VPW
MM0 ZN B net13 VPW n18 W=2.27u L=180.00n
MM13 net13 A1 VSS VPW n18 W=2.16u L=180.00n
MM12 net13 A2 VSS VPW n18 W=2.16u L=180.00n
MM2 net28 A2 VDD VNW p18 W=2.96u L=180.00n
MM1 ZN B VDD VNW p18 W=2.28u L=180.00n
MM10 ZN A1 net28 VNW p18 W=3.03u L=180.00n
.ENDS OAI21UHDV3
.SUBCKT OAI21UHDV4 A1 A2 B ZN VDD VSS VNW VPW
MM0 ZN B net13 VPW n18 W=3.11u L=180.00n
MM13 net13 A1 VSS VPW n18 W=2.88u L=180.00n
MM12 net13 A2 VSS VPW n18 W=2.88u L=180.00n
MM2 net28 A2 VDD VNW p18 W=3.88u L=180.00n
MM1 ZN B VDD VNW p18 W=2.76u L=180.00n
MM10 ZN A1 net28 VNW p18 W=4.04u L=180.00n
.ENDS OAI21UHDV4
.SUBCKT OAI21UHDV6 A1 A2 B ZN VDD VSS VNW VPW
MM0 ZN B net13 VPW n18 W=4.26u L=180.00n
MM13 net13 A1 VSS VPW n18 W=4.32u L=180.00n
MM12 net13 A2 VSS VPW n18 W=4.32u L=180.00n
MM2 net28 A2 VDD VNW p18 W=5.9u L=180.00n
MM1 ZN B VDD VNW p18 W=4.42u L=180.00n
MM10 ZN A1 net28 VNW p18 W=6.06u L=180.00n
.ENDS OAI21UHDV6
.SUBCKT OAI221UHDV0P4 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM9 net7 B2 net10 VPW n18 W=0.28u L=180.00n
MM6 net7 B1 net10 VPW n18 W=0.28u L=180.00n
MM5 ZN C net7 VPW n18 W=0.28u L=180.00n
MM4 net10 A1 VSS VPW n18 W=0.28u L=180.00n
MM3 net10 A2 VSS VPW n18 W=0.28u L=180.00n
MM8 ZN B1 net30 VNW p18 W=490.0n L=180.00n
MM2 net30 B2 VDD VNW p18 W=490.0n L=180.00n
MM1 ZN C VDD VNW p18 W=490.0n L=180.00n
MM0 ZN A1 net42 VNW p18 W=490.0n L=180.00n
MM7 net42 A2 VDD VNW p18 W=490.0n L=180.00n
.ENDS OAI221UHDV0P4
.SUBCKT OAI221UHDV0P7 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM7 net14 A2 VDD VNW p18 W=790.0n L=180.00n
MM0 ZN A1 net14 VNW p18 W=790.0n L=180.00n
MM1 ZN C VDD VNW p18 W=540.0n L=180.00n
MM2 net26 B2 VDD VNW p18 W=790.0n L=180.00n
MM8 ZN B1 net26 VNW p18 W=790.0n L=180.00n
MM5 ZN C net43 VPW n18 W=560.00n L=180.00n
MM3 net46 A2 VSS VPW n18 W=560.00n L=180.00n
MM4 net46 A1 VSS VPW n18 W=560.00n L=180.00n
MM6 net43 B1 net46 VPW n18 W=560.00n L=180.00n
MM9 net43 B2 net46 VPW n18 W=470.00n L=180.00n
.ENDS OAI221UHDV0P7
.SUBCKT OAI221UHDV1 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM7 net14 A2 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN A1 net14 VNW p18 W=1.01u L=180.00n
MM1 ZN C VDD VNW p18 W=925.00n L=180.00n
MM2 net26 B2 VDD VNW p18 W=925.00n L=180.00n
MM8 ZN B1 net26 VNW p18 W=925.00n L=180.00n
MM5 ZN C net43 VPW n18 W=720.00n L=180.00n
MM3 net46 A2 VSS VPW n18 W=720.00n L=180.00n
MM4 net46 A1 VSS VPW n18 W=720.00n L=180.00n
MM6 net43 B1 net46 VPW n18 W=0.72u L=180.00n
MM9 net43 B2 net46 VPW n18 W=770.00n L=180.00n
.ENDS OAI221UHDV1
.SUBCKT OAI221UHDV2 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM7 net14 A2 VDD VNW p18 W=1.99u L=180.00n
MM0 ZN A1 net14 VNW p18 W=1.54u L=180.00n
MM1 ZN C VDD VNW p18 W=1.85u L=180.00n
MM2 net26 B2 VDD VNW p18 W=1.74u L=180.00n
MM8 ZN B1 net26 VNW p18 W=1.85u L=180.00n
MM5 ZN C net43 VPW n18 W=1.52u L=180.00n
MM3 net46 A2 VSS VPW n18 W=1.44u L=180.00n
MM4 net46 A1 VSS VPW n18 W=1.44u L=180.00n
MM6 net43 B1 net46 VPW n18 W=1.55u L=180.00n
MM9 net43 B2 net46 VPW n18 W=1.55u L=180.00n
.ENDS OAI221UHDV2
.SUBCKT OAI221UHDV3 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM7 net14 A2 VDD VNW p18 W=3.03u L=180.00n
MM0 ZN A1 net14 VNW p18 W=2.55u L=180.00n
MM1 ZN C VDD VNW p18 W=2.775u L=180.00n
MM2 net26 B2 VDD VNW p18 W=2.335u L=180.00n
MM8 ZN B1 net26 VNW p18 W=2.77u L=180.00n
MM5 ZN C net43 VPW n18 W=2.27u L=180.00n
MM3 net46 A2 VSS VPW n18 W=2.16u L=180.00n
MM4 net46 A1 VSS VPW n18 W=2.16u L=180.00n
MM6 net43 B1 net46 VPW n18 W=2.54u L=180.00n
MM9 net43 B2 net46 VPW n18 W=2.54u L=180.00n
.ENDS OAI221UHDV3
.SUBCKT OAI221UHDV4 A1 A2 B1 B2 C ZN VDD VSS VNW VPW
MM5 ZN C net43 VPW n18 W=3u L=180.00n
MM3 net46 A2 VSS VPW n18 W=3u L=180.00n
MM4 net46 A1 VSS VPW n18 W=3u L=180.00n
MM6 net43 B1 net46 VPW n18 W=3u L=180.00n
MM9 net43 B2 net46 VPW n18 W=3u L=180.00n
MM7 net14 A2 VDD VNW p18 W=4u L=180.00n
MM0 ZN A1 net14 VNW p18 W=3.8u L=180.00n
MM1 ZN C VDD VNW p18 W=4u L=180.00n
MM2 net26 B2 VDD VNW p18 W=4u L=180.00n
MM8 ZN B1 net26 VNW p18 W=4u L=180.00n
.ENDS OAI221UHDV4
.SUBCKT OAI222UHDV0P4 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM11 ZN C1 net16 VPW n18 W=0.28u L=180.00n
MM13 net16 B1 net24 VPW n18 W=0.28u L=180.00n
MM12 net16 B2 net24 VPW n18 W=0.28u L=180.00n
MM6 ZN C2 net16 VPW n18 W=0.28u L=180.00n
MM3 net24 A2 VSS VPW n18 W=0.28u L=180.00n
MM4 net24 A1 VSS VPW n18 W=0.28u L=180.00n
MM10 ZN B1 net35 VNW p18 W=490.0n L=180.00n
MM7 net43 C2 VDD VNW p18 W=490.0n L=180.00n
MM0 ZN C1 net43 VNW p18 W=490.0n L=180.00n
MM1 net55 A2 VDD VNW p18 W=490.0n L=180.00n
MM2 net35 B2 VDD VNW p18 W=490.0n L=180.00n
MM5 ZN A1 net55 VNW p18 W=490.0n L=180.00n
.ENDS OAI222UHDV0P4
.SUBCKT OAI222UHDV0P7 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM5 ZN A1 net11 VNW p18 W=790.0n L=180.00n
MM2 net31 B2 VDD VNW p18 W=790.0n L=180.00n
MM1 net11 A2 VDD VNW p18 W=790.0n L=180.00n
MM0 ZN C1 net23 VNW p18 W=790.0n L=180.00n
MM7 net23 C2 VDD VNW p18 W=790.0n L=180.00n
MM10 ZN B1 net31 VNW p18 W=790.0n L=180.00n
MM4 net36 A1 VSS VPW n18 W=400.00n L=180.00n
MM3 net36 A2 VSS VPW n18 W=400.00n L=180.00n
MM6 ZN C2 net44 VPW n18 W=0.385u L=180.00n
MM12 net44 B2 net36 VPW n18 W=470.00n L=180.00n
MM13 net44 B1 net36 VPW n18 W=470.00n L=180.00n
MM11 ZN C1 net44 VPW n18 W=0.395u L=180.00n
.ENDS OAI222UHDV0P7
.SUBCKT OAI222UHDV1 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM5 ZN A1 net11 VNW p18 W=1.01u L=180.00n
MM2 net31 B2 VDD VNW p18 W=0.92u L=180.00n
MM1 net11 A2 VDD VNW p18 W=1.01u L=180.00n
MM0 ZN C1 net23 VNW p18 W=0.92u L=180.00n
MM7 net23 C2 VDD VNW p18 W=0.92u L=180.00n
MM10 ZN B1 net31 VNW p18 W=0.92u L=180.00n
MM4 net36 A1 VSS VPW n18 W=0.42u L=180.00n
MM3 net36 A2 VSS VPW n18 W=0.42u L=180.00n
MM6 ZN C2 net44 VPW n18 W=720.00n L=180.00n
MM12 net44 B2 net36 VPW n18 W=720.00n L=180.00n
MM13 net44 B1 net36 VPW n18 W=770.00n L=180.00n
MM11 ZN C1 net44 VPW n18 W=770.00n L=180.00n
.ENDS OAI222UHDV1
.SUBCKT OAI222UHDV2 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM5 ZN A1 net11 VNW p18 W=1.775u L=180.00n
MM2 net31 B2 VDD VNW p18 W=1.8u L=180.00n
MM1 net11 A2 VDD VNW p18 W=1.965u L=180.00n
MM0 ZN C1 net23 VNW p18 W=1.69u L=180.00n
MM7 net23 C2 VDD VNW p18 W=1.69u L=180.00n
MM10 ZN B1 net31 VNW p18 W=1.69u L=180.00n
MM4 net36 A1 VSS VPW n18 W=1.44u L=180.00n
MM3 net36 A2 VSS VPW n18 W=1.44u L=180.00n
MM6 ZN C2 net44 VPW n18 W=1.55u L=180.00n
MM12 net44 B2 net36 VPW n18 W=1.605u L=180.00n
MM13 net44 B1 net36 VPW n18 W=1.605u L=180.00n
MM11 ZN C1 net44 VPW n18 W=1.49u L=180.00n
.ENDS OAI222UHDV2
.SUBCKT OAI222UHDV3 A1 A2 B1 B2 C1 C2 ZN VDD VSS VNW VPW
MM5 ZN A1 net11 VNW p18 W=3.03u L=180.00n
MM2 net31 B2 VDD VNW p18 W=2.77u L=180.00n
MM1 net11 A2 VDD VNW p18 W=2.78u L=180.00n
MM0 ZN C1 net23 VNW p18 W=2.77u L=180.00n
MM7 net23 C2 VDD VNW p18 W=2.61u L=180.00n
MM10 ZN B1 net31 VNW p18 W=2.55u L=180.00n
MM4 net36 A1 VSS VPW n18 W=2.16u L=180.00n
MM3 net36 A2 VSS VPW n18 W=2.16u L=180.00n
MM6 ZN C2 net44 VPW n18 W=2.27u L=180.00n
MM12 net44 B2 net36 VPW n18 W=2.27u L=180.00n
MM13 net44 B1 net36 VPW n18 W=2.33u L=180.00n
MM11 ZN C1 net44 VPW n18 W=2.33u L=180.00n
.ENDS OAI222UHDV3
.SUBCKT OAI22BBUHDV0P4 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM8 net10 B2 VSS VPW n18 W=0.28u L=180.00n
MM4 net10 B1 VSS VPW n18 W=0.28u L=180.00n
MM3 ZN net42 net10 VPW n18 W=0.28u L=180.00n
MM1 net18 A2 VSS VPW n18 W=0.28u L=180.00n
MM12 net42 A1 net18 VPW n18 W=0.28u L=180.00n
MM6 ZN B1 net33 VNW p18 W=490.0n L=180.00n
MM5 ZN net42 VDD VNW p18 W=490.0n L=180.00n
MM7 net33 B2 VDD VNW p18 W=490.0n L=180.00n
MM0 net42 A2 VDD VNW p18 W=490.0n L=180.00n
MM2 net42 A1 VDD VNW p18 W=490.0n L=180.00n
.ENDS OAI22BBUHDV0P4
.SUBCKT OAI22BBUHDV0P7 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM2 net6 A1 VDD VNW p18 W=500.0n L=180.00n
MM0 net6 A2 VDD VNW p18 W=500.0n L=180.00n
MM5 ZN net6 VDD VNW p18 W=790.0n L=180.00n
MM6 ZN B1 net21 VNW p18 W=790.0n L=180.00n
MM7 net21 B2 VDD VNW p18 W=790.0n L=180.00n
MM12 net6 A1 net30 VPW n18 W=430.00n L=180.00n
MM1 net30 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 ZN net6 net38 VPW n18 W=560.00n L=180.00n
MM4 net38 B1 VSS VPW n18 W=420.00n L=180.00n
MM8 net38 B2 VSS VPW n18 W=420.00n L=180.00n
.ENDS OAI22BBUHDV0P7
.SUBCKT OAI22BBUHDV1 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM2 net6 A1 VDD VNW p18 W=580.0n L=180.00n
MM0 net6 A2 VDD VNW p18 W=580.0n L=180.00n
MM5 ZN net6 VDD VNW p18 W=1.01u L=180.00n
MM6 ZN B1 net21 VNW p18 W=1.01u L=180.00n
MM7 net21 B2 VDD VNW p18 W=1.01u L=180.00n
MM12 net6 A1 net30 VPW n18 W=430.00n L=180.00n
MM1 net30 A2 VSS VPW n18 W=430.00n L=180.00n
MM3 ZN net6 net38 VPW n18 W=720.00n L=180.00n
MM4 net38 B1 VSS VPW n18 W=720.00n L=180.00n
MM8 net38 B2 VSS VPW n18 W=720.00n L=180.00n
.ENDS OAI22BBUHDV1
.SUBCKT OAI22BBUHDV2 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM2 net6 A1 VDD VNW p18 W=950.0n L=180.00n
MM0 net6 A2 VDD VNW p18 W=950.0n L=180.00n
MM5 ZN net6 VDD VNW p18 W=1.9u L=180.00n
MM6 ZN B1 net21 VNW p18 W=2.02u L=180.00n
MM7 net21 B2 VDD VNW p18 W=1.985u L=180.00n
MM12 net6 A1 net30 VPW n18 W=630.00n L=180.00n
MM1 net30 A2 VSS VPW n18 W=630.00n L=180.00n
MM3 ZN net6 net38 VPW n18 W=1.55u L=180.00n
MM4 net38 B1 VSS VPW n18 W=1.39u L=180.00n
MM8 net38 B2 VSS VPW n18 W=1.415u L=180.00n
.ENDS OAI22BBUHDV2
.SUBCKT OAI22UHDV0P4 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM5 ZN A1 net9 VNW p18 W=490.0n L=180.00n
MM2 net21 B2 VDD VNW p18 W=490.0n L=180.00n
MM1 net9 A2 VDD VNW p18 W=490.0n L=180.00n
MM10 ZN B1 net21 VNW p18 W=490.0n L=180.00n
MM11 ZN B1 net30 VPW n18 W=0.28u L=180.00n
MM6 ZN B2 net30 VPW n18 W=0.25u L=180.00n
MM12 net30 A2 VSS VPW n18 W=0.28u L=180.00n
MM13 net30 A1 VSS VPW n18 W=0.28u L=180.00n
.ENDS OAI22UHDV0P4
.SUBCKT OAI22UHDV0P7 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM13 net10 A1 VSS VPW n18 W=560.00n L=180.00n
MM12 net10 A2 VSS VPW n18 W=560.00n L=180.00n
MM6 ZN B2 net10 VPW n18 W=560.00n L=180.00n
MM11 ZN B1 net10 VPW n18 W=560.00n L=180.00n
MM10 ZN B1 net25 VNW p18 W=790.0n L=180.00n
MM1 net37 A2 VDD VNW p18 W=790.0n L=180.00n
MM2 net25 B2 VDD VNW p18 W=790.0n L=180.00n
MM5 ZN A1 net37 VNW p18 W=790.0n L=180.00n
.ENDS OAI22UHDV0P7
.SUBCKT OAI22UHDV1 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM13 net10 A1 VSS VPW n18 W=720.00n L=180.00n
MM12 net10 A2 VSS VPW n18 W=720.00n L=180.00n
MM6 ZN B2 net10 VPW n18 W=0.72u L=180.00n
MM11 ZN B1 net10 VPW n18 W=0.72u L=180.00n
MM10 ZN B1 net25 VNW p18 W=0.92u L=180.00n
MM1 net37 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net25 B2 VDD VNW p18 W=0.92u L=180.00n
MM5 ZN A1 net37 VNW p18 W=1.01u L=180.00n
.ENDS OAI22UHDV1
.SUBCKT OAI22UHDV2 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM13 net10 A1 VSS VPW n18 W=1.44u L=180.00n
MM12 net10 A2 VSS VPW n18 W=1.44u L=180.00n
MM6 ZN B2 net10 VPW n18 W=1.5u L=180.00n
MM11 ZN B1 net10 VPW n18 W=1.55u L=180.00n
MM10 ZN B1 net25 VNW p18 W=1.53u L=180.00n
MM1 net37 A2 VDD VNW p18 W=1.94u L=180.00n
MM2 net25 B2 VDD VNW p18 W=1.685u L=180.00n
MM5 ZN A1 net37 VNW p18 W=1.94u L=180.00n
.ENDS OAI22UHDV2
.SUBCKT OAI22UHDV3 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM13 net10 A1 VSS VPW n18 W=2.16u L=180.00n
MM12 net10 A2 VSS VPW n18 W=2.16u L=180.00n
MM6 ZN B2 net10 VPW n18 W=2.16u L=180.00n
MM11 ZN B1 net10 VPW n18 W=2.16u L=180.00n
MM10 ZN B1 net25 VNW p18 W=2.45u L=180.00n
MM1 net37 A2 VDD VNW p18 W=2.51u L=180.00n
MM2 net25 B2 VDD VNW p18 W=2.76u L=180.00n
MM5 ZN A1 net37 VNW p18 W=2.9u L=180.00n
.ENDS OAI22UHDV3
.SUBCKT OAI22UHDV4 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM13 net10 A1 VSS VPW n18 W=2.88u L=180.00n
MM12 net10 A2 VSS VPW n18 W=2.88u L=180.00n
MM6 ZN B2 net10 VPW n18 W=3.11u L=180.00n
MM11 ZN B1 net10 VPW n18 W=3.11u L=180.00n
MM10 ZN B1 net25 VNW p18 W=3.06u L=180.00n
MM1 net37 A2 VDD VNW p18 W=3.955u L=180.00n
MM2 net25 B2 VDD VNW p18 W=3.7u L=180.00n
MM5 ZN A1 net37 VNW p18 W=3.48u L=180.00n
.ENDS OAI22UHDV4
.SUBCKT OAI22UHDV6 A1 A2 B1 B2 ZN VDD VSS VNW VPW
MM13 net10 A1 VSS VPW n18 W=4.32u L=180.00n
MM12 net10 A2 VSS VPW n18 W=4.32u L=180.00n
MM6 ZN B2 net10 VPW n18 W=4.66u L=180.00n
MM11 ZN B1 net10 VPW n18 W=4.66u L=180.00n
MM10 ZN B1 net25 VNW p18 W=4.59u L=180.00n
MM1 net37 A2 VDD VNW p18 W=5.835u L=180.00n
MM2 net25 B2 VDD VNW p18 W=5.55u L=180.00n
MM5 ZN A1 net37 VNW p18 W=5.22u L=180.00n
.ENDS OAI22UHDV6
.SUBCKT OAI22XBUHDV0P4 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM3 B2 B2N VSS VPW n18 W=250.00n L=180.00n
MM13 net10 A1 VSS VPW n18 W=290.00n L=180.00n
MM12 net10 A2 VSS VPW n18 W=290.00n L=180.00n
MM6 ZN B2 net10 VPW n18 W=290.00n L=180.00n
MM11 ZN B1 net10 VPW n18 W=290.00n L=180.00n
MM0 B2 B2N VDD VNW p18 W=250.00n L=180.00n
MM10 ZN B1 net25 VNW p18 W=400.00n L=180.00n
MM1 net37 A2 VDD VNW p18 W=400.00n L=180.00n
MM2 net25 B2 VDD VNW p18 W=400.00n L=180.00n
MM5 ZN A1 net37 VNW p18 W=400.00n L=180.00n
.ENDS OAI22XBUHDV0P4
.SUBCKT OAI22XBUHDV0P7 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM3 B2 B2N VSS VPW n18 W=250.00n L=180.00n
MM13 net10 A1 VSS VPW n18 W=500.00n L=180.00n
MM12 net10 A2 VSS VPW n18 W=500.00n L=180.00n
MM6 ZN B2 net10 VPW n18 W=500.00n L=180.00n
MM11 ZN B1 net10 VPW n18 W=500.00n L=180.00n
MM0 B2 B2N VDD VNW p18 W=280.00n L=180.00n
MM10 ZN B1 net25 VNW p18 W=710.00n L=180.00n
MM1 net37 A2 VDD VNW p18 W=710.00n L=180.00n
MM2 net25 B2 VDD VNW p18 W=710.00n L=180.00n
MM5 ZN A1 net37 VNW p18 W=710.00n L=180.00n
.ENDS OAI22XBUHDV0P7
.SUBCKT OAI22XBUHDV1 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM3 B2 B2N VSS VPW n18 W=290.00n L=180.00n
MM13 net10 A1 VSS VPW n18 W=720.00n L=180.00n
MM12 net10 A2 VSS VPW n18 W=720.00n L=180.00n
MM6 ZN B2 net10 VPW n18 W=720.00n L=180.00n
MM11 ZN B1 net10 VPW n18 W=720.00n L=180.00n
MM0 B2 B2N VDD VNW p18 W=410.00n L=180.00n
MM10 ZN B1 net25 VNW p18 W=0.95u L=180.00n
MM1 net37 A2 VDD VNW p18 W=1.01u L=180.00n
MM2 net25 B2 VDD VNW p18 W=0.95u L=180.00n
MM5 ZN A1 net37 VNW p18 W=0.95u L=180.00n
.ENDS OAI22XBUHDV1
.SUBCKT OAI22XBUHDV2 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM3 B2 B2N VSS VPW n18 W=580.00n L=180.00n
MM13 net10 A1 VSS VPW n18 W=1.44u L=180.00n
MM12 net10 A2 VSS VPW n18 W=1.44u L=180.00n
MM6 ZN B2 net10 VPW n18 W=1.44u L=180.00n
MM11 ZN B1 net10 VPW n18 W=1.44u L=180.00n
MM0 B2 B2N VDD VNW p18 W=810.00n L=180.00n
MM10 ZN B1 net25 VNW p18 W=1.86u L=180.00n
MM1 net37 A2 VDD VNW p18 W=1.95u L=180.00n
MM2 net25 B2 VDD VNW p18 W=1.86u L=180.00n
MM5 ZN A1 net37 VNW p18 W=1.95u L=180.00n
.ENDS OAI22XBUHDV2
.SUBCKT OAI22XBUHDV4 A1 A2 B1 B2N ZN VDD VSS VNW VPW
MM3 B2 B2N VSS VPW n18 W=1.16u L=180.00n
MM13 net10 A1 VSS VPW n18 W=2.88u L=180.00n
MM12 net10 A2 VSS VPW n18 W=2.88u L=180.00n
MM6 ZN B2 net10 VPW n18 W=2.88u L=180.00n
MM11 ZN B1 net10 VPW n18 W=2.88u L=180.00n
MM0 B2 B2N VDD VNW p18 W=1.62u L=180.00n
MM10 ZN B1 net25 VNW p18 W=3.08u L=180.00n
MM1 net37 A2 VDD VNW p18 W=3.9u L=180.00n
MM2 net25 B2 VDD VNW p18 W=3.72u L=180.00n
MM5 ZN A1 net37 VNW p18 W=3.9u L=180.00n
.ENDS OAI22XBUHDV4
.SUBCKT OAI2XB11UHDV0P4 A1 A2N B C ZN VDD VSS VNW VPW
MM8 net063 A2N VSS VPW n18 W=250.00n L=180.00n
MM6 net6 B net18 VPW n18 W=290.00n L=180.00n
MM5 ZN C net6 VPW n18 W=290.00n L=180.00n
MM4 net18 A1 VSS VPW n18 W=290.00n L=180.00n
MM3 net18 net063 VSS VPW n18 W=290.00n L=180.00n
MM9 net063 A2N VDD VNW p18 W=250.00n L=180.00n
MM2 ZN C VDD VNW p18 W=400.00n L=180.00n
MM1 ZN B VDD VNW p18 W=400.00n L=180.00n
MM0 ZN A1 net33 VNW p18 W=400.00n L=180.00n
MM7 net33 net063 VDD VNW p18 W=400.00n L=180.00n
.ENDS OAI2XB11UHDV0P4
.SUBCKT OAI2XB11UHDV0P7 A1 A2N B C ZN VDD VSS VNW VPW
MM8 net063 A2N VSS VPW n18 W=250.00n L=180.00n
MM6 net6 B net18 VPW n18 W=500.00n L=180.00n
MM5 ZN C net6 VPW n18 W=500.00n L=180.00n
MM4 net18 A1 VSS VPW n18 W=500.00n L=180.00n
MM3 net18 net063 VSS VPW n18 W=500.00n L=180.00n
MM9 net063 A2N VDD VNW p18 W=280.00n L=180.00n
MM2 ZN C VDD VNW p18 W=710.00n L=180.00n
MM1 ZN B VDD VNW p18 W=710.00n L=180.00n
MM0 ZN A1 net33 VNW p18 W=710.00n L=180.00n
MM7 net33 net063 VDD VNW p18 W=710.00n L=180.00n
.ENDS OAI2XB11UHDV0P7
.SUBCKT OAI2XB11UHDV1 A1 A2N B C ZN VDD VSS VNW VPW
MM8 net063 A2N VSS VPW n18 W=290.00n L=180.00n
MM6 net6 B net18 VPW n18 W=720.00n L=180.00n
MM5 ZN C net6 VPW n18 W=720.00n L=180.00n
MM4 net18 A1 VSS VPW n18 W=720.00n L=180.00n
MM3 net18 net063 VSS VPW n18 W=720.00n L=180.00n
MM9 net063 A2N VDD VNW p18 W=410.00n L=180.00n
MM2 ZN C VDD VNW p18 W=1.01u L=180.00n
MM1 ZN B VDD VNW p18 W=1.01u L=180.00n
MM0 ZN A1 net33 VNW p18 W=1.01u L=180.00n
MM7 net33 net063 VDD VNW p18 W=1.01u L=180.00n
.ENDS OAI2XB11UHDV1
.SUBCKT OAI2XB11UHDV2 A1 A2N B C ZN VDD VSS VNW VPW
MM8 net063 A2N VSS VPW n18 W=580.00n L=180.00n
MM6 net6 B net18 VPW n18 W=1.44u L=180.00n
MM5 ZN C net6 VPW n18 W=1.44u L=180.00n
MM4 net18 A1 VSS VPW n18 W=1.44u L=180.00n
MM3 net18 net063 VSS VPW n18 W=1.44u L=180.00n
MM9 net063 A2N VDD VNW p18 W=810.00n L=180.00n
MM2 ZN C VDD VNW p18 W=1.9u L=180.00n
MM1 ZN B VDD VNW p18 W=2.02u L=180.00n
MM0 ZN A1 net33 VNW p18 W=2.02u L=180.00n
MM7 net33 net063 VDD VNW p18 W=2.02u L=180.00n
.ENDS OAI2XB11UHDV2
.SUBCKT OAI2XB1UHDV0P4 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VSS VPW n18 W=250.00n L=180.00n
MM0 ZN A net13 VPW n18 W=290.00n L=180.00n
MM13 net13 B1 VSS VPW n18 W=290.00n L=180.00n
MM12 net13 b2n VSS VPW n18 W=290.00n L=180.00n
MM3 b2n B2 VDD VNW p18 W=250.00n L=180.00n
MM2 net28 b2n VDD VNW p18 W=400.00n L=180.00n
MM1 ZN A VDD VNW p18 W=400.00n L=180.00n
MM10 ZN B1 net28 VNW p18 W=400.00n L=180.00n
.ENDS OAI2XB1UHDV0P4
.SUBCKT OAI2XB1UHDV0P7 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VSS VPW n18 W=250.00n L=180.00n
MM0 ZN A net13 VPW n18 W=500.00n L=180.00n
MM13 net13 B1 VSS VPW n18 W=500.00n L=180.00n
MM12 net13 b2n VSS VPW n18 W=500.00n L=180.00n
MM3 b2n B2 VDD VNW p18 W=280.00n L=180.00n
MM2 net28 b2n VDD VNW p18 W=710.00n L=180.00n
MM1 ZN A VDD VNW p18 W=710.00n L=180.00n
MM10 ZN B1 net28 VNW p18 W=710.00n L=180.00n
.ENDS OAI2XB1UHDV0P7
.SUBCKT OAI2XB1UHDV1 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VSS VPW n18 W=290.00n L=180.00n
MM0 ZN A net13 VPW n18 W=720.00n L=180.00n
MM13 net13 B1 VSS VPW n18 W=720.00n L=180.00n
MM12 net13 b2n VSS VPW n18 W=720.00n L=180.00n
MM3 b2n B2 VDD VNW p18 W=410.00n L=180.00n
MM2 net28 b2n VDD VNW p18 W=1.01u L=180.00n
MM1 ZN A VDD VNW p18 W=1.01u L=180.00n
MM10 ZN B1 net28 VNW p18 W=1.01u L=180.00n
.ENDS OAI2XB1UHDV1
.SUBCKT OAI2XB1UHDV2 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VSS VPW n18 W=580.00n L=180.00n
MM0 ZN A net13 VPW n18 W=1.44u L=180.00n
MM13 net13 B1 VSS VPW n18 W=1.44u L=180.00n
MM12 net13 b2n VSS VPW n18 W=1.44u L=180.00n
MM3 b2n B2 VDD VNW p18 W=810.00n L=180.00n
MM2 net28 b2n VDD VNW p18 W=2.02u L=180.00n
MM1 ZN A VDD VNW p18 W=1.9u L=180.00n
MM10 ZN B1 net28 VNW p18 W=2.02u L=180.00n
.ENDS OAI2XB1UHDV2
.SUBCKT OAI2XB1UHDV4 A B1 B2 ZN VDD VSS VNW VPW
MM4 b2n B2 VSS VPW n18 W=1.16u L=180.00n
MM0 ZN A net13 VPW n18 W=3.23u L=180.00n
MM13 net13 B1 VSS VPW n18 W=2.88u L=180.00n
MM12 net13 b2n VSS VPW n18 W=2.88u L=180.00n
MM3 b2n B2 VDD VNW p18 W=1.62u L=180.00n
MM2 net28 b2n VDD VNW p18 W=3.97u L=180.00n
MM1 ZN A VDD VNW p18 W=3.72u L=180.00n
MM10 ZN B1 net28 VNW p18 W=3.97u L=180.00n
.ENDS OAI2XB1UHDV4
.SUBCKT OAI31UHDV0P4 A1 A2 A3 B ZN VDD VSS VNW VPW
MM4 net6 A3 VSS VPW n18 W=0.265u L=180.00n
MM0 ZN B net6 VPW n18 W=0.28u L=180.00n
MM13 net6 A1 VSS VPW n18 W=0.42u L=180.00n
MM12 net6 A2 VSS VPW n18 W=0.28u L=180.00n
MM3 net33 A3 VDD VNW p18 W=490.0n L=180.00n
MM2 net37 A2 net33 VNW p18 W=490.0n L=180.00n
MM1 ZN B VDD VNW p18 W=490.0n L=180.00n
MM10 ZN A1 net37 VNW p18 W=490.0n L=180.00n
.ENDS OAI31UHDV0P4
.SUBCKT OAI31UHDV0P7 A1 A2 A3 B ZN VDD VSS VNW VPW
MM10 ZN A1 net9 VNW p18 W=790.0n L=180.00n
MM2 net9 A2 net13 VNW p18 W=790.0n L=180.00n
MM3 net13 A3 VDD VNW p18 W=790.0n L=180.00n
MM1 ZN B VDD VNW p18 W=790.00n L=180.00n
MM0 ZN B net34 VPW n18 W=560.00n L=180.00n
MM12 net34 A2 VSS VPW n18 W=0.56u L=180.00n
MM13 net34 A1 VSS VPW n18 W=0.56u L=180.00n
MM4 net34 A3 VSS VPW n18 W=560.00n L=180.00n
.ENDS OAI31UHDV0P7
.SUBCKT OAI31UHDV1 A1 A2 A3 B ZN VDD VSS VNW VPW
MM10 ZN A1 net9 VNW p18 W=1.01u L=180.00n
MM2 net9 A2 net13 VNW p18 W=1.01u L=180.00n
MM3 net13 A3 VDD VNW p18 W=1.01u L=180.00n
MM1 ZN B VDD VNW p18 W=1.01u L=180.00n
MM0 ZN B net34 VPW n18 W=720.00n L=180.00n
MM12 net34 A2 VSS VPW n18 W=720.00n L=180.00n
MM13 net34 A1 VSS VPW n18 W=720.00n L=180.00n
MM4 net34 A3 VSS VPW n18 W=720.00n L=180.00n
.ENDS OAI31UHDV1
.SUBCKT OAI31UHDV2 A1 A2 A3 B ZN VDD VSS VNW VPW
MM10 ZN A1 net9 VNW p18 W=1.52u L=180.00n
MM2 net9 A2 net13 VNW p18 W=1.89u L=180.00n
MM3 net13 A3 VDD VNW p18 W=1.93u L=180.00n
MM1 ZN B VDD VNW p18 W=1.85u L=180.00n
MM0 ZN B net34 VPW n18 W=1.55u L=180.00n
MM12 net34 A2 VSS VPW n18 W=1.44u L=180.00n
MM13 net34 A1 VSS VPW n18 W=1.44u L=180.00n
MM4 net34 A3 VSS VPW n18 W=1.44u L=180.00n
.ENDS OAI31UHDV2
.SUBCKT OAI31UHDV3 A1 A2 A3 B ZN VDD VSS VNW VPW
MM10 ZN A1 net9 VNW p18 W=3.03u L=180.00n
MM2 net9 A2 net13 VNW p18 W=3.03u L=180.00n
MM3 net13 A3 VDD VNW p18 W=3.03u L=180.00n
MM1 ZN B VDD VNW p18 W=2.775u L=180.00n
MM0 ZN B net34 VPW n18 W=2.27u L=180.00n
MM12 net34 A2 VSS VPW n18 W=2.16u L=180.00n
MM13 net34 A1 VSS VPW n18 W=2.16u L=180.00n
MM4 net34 A3 VSS VPW n18 W=2.16u L=180.00n
.ENDS OAI31UHDV3
****Sub-Circuit for OAI32UHDV0P4, Tue Jun  6 16:00:22 CST 2017****
.SUBCKT OAI32UHDV0P4 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM6 ZN B1 net34 VPW n18 W=290.00n L=180.00n
MM0 ZN B2 net34 VPW n18 W=290.00n L=180.00n
MM12 net34 A2 VSS VPW n18 W=290.00n L=180.00n
MM13 net34 A1 VSS VPW n18 W=290.00n L=180.00n
MM4 net34 A3 VSS VPW n18 W=290.00n L=180.00n
MM5 ZN B1 net040 VNW p18 W=490.00n L=180.00n
MM10 ZN A1 net9 VNW p18 W=490.00n L=180.00n
MM2 net9 A2 net13 VNW p18 W=490.00n L=180.00n
MM3 net13 A3 VDD VNW p18 W=490.00n L=180.00n
MM1 net040 B2 VDD VNW p18 W=490.00n L=180.00n
.ENDS OAI32UHDV0P4
****Sub-Circuit for OAI32UHDV0P7, Tue Jun  6 16:00:22 CST 2017****
.SUBCKT OAI32UHDV0P7 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM6 ZN B1 net34 VPW n18 W=560.00n L=180.00n
MM0 ZN B2 net34 VPW n18 W=560.00n L=180.00n
MM12 net34 A2 VSS VPW n18 W=560.00n L=180.00n
MM13 net34 A1 VSS VPW n18 W=560.00n L=180.00n
MM4 net34 A3 VSS VPW n18 W=560.00n L=180.00n
MM5 ZN B1 net040 VNW p18 W=790.00n L=180.00n
MM10 ZN A1 net9 VNW p18 W=790.00n L=180.00n
MM2 net9 A2 net13 VNW p18 W=790.00n L=180.00n
MM3 net13 A3 VDD VNW p18 W=790.00n L=180.00n
MM1 net040 B2 VDD VNW p18 W=790.00n L=180.00n
.ENDS OAI32UHDV0P7
****Sub-Circuit for OAI32UHDV1, Tue Jun  6 16:00:22 CST 2017****
.SUBCKT OAI32UHDV1 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM6 ZN B1 net34 VPW n18 W=720.00n L=180.00n
MM0 ZN B2 net34 VPW n18 W=720.00n L=180.00n
MM12 net34 A2 VSS VPW n18 W=720.00n L=180.00n
MM13 net34 A1 VSS VPW n18 W=720.00n L=180.00n
MM4 net34 A3 VSS VPW n18 W=720.00n L=180.00n
MM5 ZN B1 net040 VNW p18 W=950.00n L=180.00n
MM10 ZN A1 net9 VNW p18 W=1.01u L=180.00n
MM2 net9 A2 net13 VNW p18 W=1.01u L=180.00n
MM3 net13 A3 VDD VNW p18 W=1.01u L=180.00n
MM1 net040 B2 VDD VNW p18 W=950.00n L=180.00n
.ENDS OAI32UHDV1
****Sub-Circuit for OAI32UHDV2, Tue Jun  6 16:00:22 CST 2017****
.SUBCKT OAI32UHDV2 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM6 ZN B1 net34 VPW n18 W=1.44u L=180.00n
MM0 ZN B2 net34 VPW n18 W=1.44u L=180.00n
MM12 net34 A2 VSS VPW n18 W=1.44u L=180.00n
MM13 net34 A1 VSS VPW n18 W=1.44u L=180.00n
MM4 net34 A3 VSS VPW n18 W=1.44u L=180.00n
MM5 ZN B1 net040 VNW p18 W=1.72u L=180.00n
MM10 ZN A1 net9 VNW p18 W=1.48u L=180.00n
MM2 net9 A2 net13 VNW p18 W=1.94u L=180.00n
MM3 net13 A3 VDD VNW p18 W=1.98u L=180.00n
MM1 net040 B2 VDD VNW p18 W=1.9u L=180.00n
.ENDS OAI32UHDV2
****Sub-Circuit for OAI32UHDV3, Tue Jun  6 16:00:22 CST 2017****
.SUBCKT OAI32UHDV3 A1 A2 A3 B1 B2 ZN VDD VSS VNW VPW
MM6 ZN B1 net34 VPW n18 W=2.16u L=180.00n
MM0 ZN B2 net34 VPW n18 W=2.16u L=180.00n
MM12 net34 A2 VSS VPW n18 W=2.16u L=180.00n
MM13 net34 A1 VSS VPW n18 W=2.16u L=180.00n
MM4 net34 A3 VSS VPW n18 W=2.16u L=180.00n
MM5 ZN B1 net040 VNW p18 W=2.85u L=180.00n
MM10 ZN A1 net9 VNW p18 W=3.03u L=180.00n
MM2 net9 A2 net13 VNW p18 W=3.03u L=180.00n
MM3 net13 A3 VDD VNW p18 W=3.03u L=180.00n
MM1 net040 B2 VDD VNW p18 W=2.85u L=180.00n
.ENDS OAI32UHDV3
.SUBCKT OR2UHDV0P4 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=0.28u L=180.00n
MM15 net8 A2 VSS VPW n18 W=0.28u L=180.00n
MM8 Z net8 VSS VPW n18 W=0.28u L=180.00n
MM0 net8 A1 net19 VNW p18 W=0.46u L=180.00n
MM7 net19 A2 VDD VNW p18 W=0.46u L=180.00n
MM6 Z net8 VDD VNW p18 W=490.00n L=180.00n
.ENDS OR2UHDV0P4
.SUBCKT OR2UHDV0P7 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=0.42u L=180.00n
MM15 net8 A2 VSS VPW n18 W=0.42u L=180.00n
MM8 Z net8 VSS VPW n18 W=560.00n L=180.00n
MM0 net8 A1 net19 VNW p18 W=500.00n L=180.00n
MM7 net19 A2 VDD VNW p18 W=500.00n L=180.00n
MM6 Z net8 VDD VNW p18 W=790.00n L=180.00n
.ENDS OR2UHDV0P7
.SUBCKT OR2UHDV1 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=0.42u L=180.00n
MM15 net8 A2 VSS VPW n18 W=0.42u L=180.00n
MM8 Z net8 VSS VPW n18 W=720.0n L=180.00n
MM0 net8 A1 net19 VNW p18 W=580.00n L=180.00n
MM7 net19 A2 VDD VNW p18 W=580.00n L=180.00n
MM6 Z net8 VDD VNW p18 W=1.01u L=180.00n
.ENDS OR2UHDV1
.SUBCKT OR2UHDV2 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=630.00n L=180.00n
MM15 net8 A2 VSS VPW n18 W=630.00n L=180.00n
MM8 Z net8 VSS VPW n18 W=1.44u L=180.00n
MM0 net8 A1 net19 VNW p18 W=0.87u L=180.00n
MM7 net19 A2 VDD VNW p18 W=0.87u L=180.00n
MM6 Z net8 VDD VNW p18 W=2.02u L=180.00n
.ENDS OR2UHDV2
.SUBCKT OR2UHDV3 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=720.00n L=180.00n
MM15 net8 A2 VSS VPW n18 W=720.00n L=180.00n
MM8 Z net8 VSS VPW n18 W=2.16u L=180.00n
MM0 net8 A1 net19 VNW p18 W=1.01u L=180.00n
MM7 net19 A2 VDD VNW p18 W=1.01u L=180.00n
MM6 Z net8 VDD VNW p18 W=3.03u L=180.00n
.ENDS OR2UHDV3
.SUBCKT OR2UHDV4 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=1.08u L=180.00n
MM15 net8 A2 VSS VPW n18 W=1.08u L=180.00n
MM8 Z net8 VSS VPW n18 W=3.2u L=180.00n
MM0 net8 A1 net19 VNW p18 W=1.49u L=180.00n
MM7 net19 A2 VDD VNW p18 W=1.49u L=180.00n
MM6 Z net8 VDD VNW p18 W=4.04u L=180.00n
.ENDS OR2UHDV4
.SUBCKT OR2UHDV6 A1 A2 Z VDD VSS VNW VPW
MM3 net8 A1 VSS VPW n18 W=1.44u L=180.00n
MM15 net8 A2 VSS VPW n18 W=1.44u L=180.00n
MM8 Z net8 VSS VPW n18 W=4.32u L=180.00n
MM0 net8 A1 net19 VNW p18 W=1.78u L=180.00n
MM7 net19 A2 VDD VNW p18 W=1.78u L=180.00n
MM6 Z net8 VDD VNW p18 W=6.06u L=180.00n
.ENDS OR2UHDV6
.SUBCKT OR2UHDV8 A1 A2 Z VDD VSS VNW VPW
MM7 net15 A2 VDD VNW p18 W=2.96u L=180.00n
MM0 net20 A1 net15 VNW p18 W=3.03u L=180.00n
MM6 Z net20 VDD VNW p18 W=8.08u L=180.00n
MM8 Z net20 VSS VPW n18 W=5.76u L=180.00n
MM15 net20 A2 VSS VPW n18 W=2.16u L=180.00n
MM3 net20 A1 VSS VPW n18 W=2.16u L=180.00n
.ENDS OR2UHDV8
.SUBCKT OR3UHDV0P7 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net12 A3 VDD VNW p18 W=500.00n L=180.00n
MM0 net16 A2 net12 VNW p18 W=500.00n L=180.00n
MM2 net21 A1 net16 VNW p18 W=500.00n L=180.00n
MM6 Z net21 VDD VNW p18 W=790.00n L=180.00n
MM15 net21 A3 VSS VPW n18 W=0.42u L=180.00n
MM3 net21 A2 VSS VPW n18 W=0.42u L=180.00n
MM4 net21 A1 VSS VPW n18 W=0.42u L=180.00n
MM8 Z net21 VSS VPW n18 W=560.00n L=180.00n
.ENDS OR3UHDV0P7
.SUBCKT OR3UHDV1 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net12 A3 VDD VNW p18 W=580.00n L=180.00n
MM0 net16 A2 net12 VNW p18 W=580.00n L=180.00n
MM2 net21 A1 net16 VNW p18 W=580.00n L=180.00n
MM6 Z net21 VDD VNW p18 W=1.01u L=180.00n
MM15 net21 A3 VSS VPW n18 W=0.42u L=180.00n
MM3 net21 A2 VSS VPW n18 W=0.42u L=180.00n
MM4 net21 A1 VSS VPW n18 W=0.42u L=180.00n
MM8 Z net21 VSS VPW n18 W=720.0n L=180.00n
.ENDS OR3UHDV1
.SUBCKT OR3UHDV2 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net12 A3 VDD VNW p18 W=0.87u L=180.00n
MM0 net16 A2 net12 VNW p18 W=0.87u L=180.00n
MM2 net21 A1 net16 VNW p18 W=0.87u L=180.00n
MM6 Z net21 VDD VNW p18 W=2.02u L=180.00n
MM15 net21 A3 VSS VPW n18 W=630.00n L=180.00n
MM3 net21 A2 VSS VPW n18 W=630.00n L=180.00n
MM4 net21 A1 VSS VPW n18 W=630.00n L=180.00n
MM8 Z net21 VSS VPW n18 W=1.44u L=180.00n
.ENDS OR3UHDV2
.SUBCKT OR3UHDV3 A1 A2 A3 Z VDD VSS VNW VPW
MM7 net12 A3 VDD VNW p18 W=1.01u L=180.00n
MM0 net16 A2 net12 VNW p18 W=1.01u L=180.00n
MM2 net21 A1 net16 VNW p18 W=1.01u L=180.00n
MM6 Z net21 VDD VNW p18 W=3.03u L=180.00n
MM15 net21 A3 VSS VPW n18 W=720.00n L=180.00n
MM3 net21 A2 VSS VPW n18 W=720.00n L=180.00n
MM4 net21 A1 VSS VPW n18 W=720.00n L=180.00n
MM8 Z net21 VSS VPW n18 W=2.16u L=180.00n
.ENDS OR3UHDV3
.SUBCKT OR3UHDV4 A1 A2 A3 Z VDD VSS VNW VPW
MM4 net17 A1 VSS VPW n18 W=1000.00n L=180.00n
MM3 net17 A2 VSS VPW n18 W=1000.00n L=180.00n
MM15 net17 A3 VSS VPW n18 W=1000.00n L=180.00n
MM8 Z net17 VSS VPW n18 W=2.88u L=180.00n
MM6 Z net17 VDD VNW p18 W=4.04u L=180.00n
MM2 net17 A1 net28 VNW p18 W=1.33u L=180.00n
MM0 net28 A2 net32 VNW p18 W=1.33u L=180.00n
MM7 net32 A3 VDD VNW p18 W=1.33u L=180.00n
.ENDS OR3UHDV4
.SUBCKT OR4UHDV0P7 A1 A2 A3 A4 Z VDD VSS VNW VPW
MM6 Z net38 VDD VNW p18 W=790.00n L=180.00n
MM2 net17 A2 net13 VNW p18 W=500.00n L=180.00n
MM1 net38 A1 net17 VNW p18 W=500.00n L=180.00n
MM0 net13 A3 net21 VNW p18 W=500.00n L=180.00n
MM7 net21 A4 VDD VNW p18 W=500.00n L=180.00n
MM5 net38 A1 VSS VPW n18 W=0.42u L=180.00n
MM4 net38 A2 VSS VPW n18 W=0.42u L=180.00n
MM3 net38 A3 VSS VPW n18 W=0.42u L=180.00n
MM15 net38 A4 VSS VPW n18 W=0.42u L=180.00n
MM8 Z net38 VSS VPW n18 W=560.00n L=180.00n
.ENDS OR4UHDV0P7
.SUBCKT OR4UHDV1 A1 A2 A3 A4 Z VDD VSS VNW VPW
MM8 Z net071 VSS VPW n18 W=720.00n L=180.00n
MM15 net071 A4 VSS VPW n18 W=0.42u L=180.00n
MM3 net071 A3 VSS VPW n18 W=0.42u L=180.00n
MM4 net071 A2 VSS VPW n18 W=0.42u L=180.00n
MM5 net071 A1 VSS VPW n18 W=0.42u L=180.00n
MM7 net29 A4 VDD VNW p18 W=580.00n L=180.00n
MM0 net37 A3 net29 VNW p18 W=580.00n L=180.00n
MM1 net071 A1 net33 VNW p18 W=580.00n L=180.00n
MM2 net33 A2 net37 VNW p18 W=580.00n L=180.00n
MM6 Z net071 VDD VNW p18 W=1.01u L=180.00n
.ENDS OR4UHDV1
.SUBCKT OR4UHDV2 A1 A2 A3 A4 Z VDD VSS VNW VPW
MM7 net54 A4 VDD VNW p18 W=0.87u L=180.00n
MM0 net46 A3 net54 VNW p18 W=0.87u L=180.00n
MM1 net71 A1 net50 VNW p18 W=0.87u L=180.00n
MM2 net50 A2 net46 VNW p18 W=0.87u L=180.00n
MM6 Z net71 VDD VNW p18 W=2.02u L=180.00n
MM8 Z net71 VSS VPW n18 W=1.44u L=180.00n
MM15 net71 A4 VSS VPW n18 W=720.00n L=180.00n
MM3 net71 A3 VSS VPW n18 W=720.00n L=180.00n
MM4 net71 A2 VSS VPW n18 W=720.00n L=180.00n
MM5 net71 A1 VSS VPW n18 W=720.00n L=180.00n
.ENDS OR4UHDV2
.SUBCKT PULLUHD0 Z VDD VSS VNW VPW
MM2 net4 net4 VDD VNW p18 W=0.42u L=180.00n
MM3 Z net4 VSS VPW n18 W=430.00n L=180.00n
.ENDS PULLUHD0
.SUBCKT PULLUHD1 Z VDD VSS VNW VPW
MM3 net4 net4 VSS VPW n18 W=430.00n L=180.00n
MM2 Z net4 VDD VNW p18 W=490.0n L=180.00n
.ENDS PULLUHD1
****Sub-Circuit for SDGRNQNUHDV0P7, Mon Jun 26 14:40:26 CST 2017****
.SUBCKT SDGRNQNUHDV0P7 CK D QN RN SE SI VDD VSS VNW VPW
MM34 net0132 RN VSS VPW n18 W=0.565u L=180.00n
MM6 net14 SEN net0132 VPW n18 W=0.565u L=180.00n
MM4 net18 cn net30 VPW n18 W=430.00n L=180.00n
MM5 net22 SI VSS VPW n18 W=430.00n L=180.00n
MM8 net30 SE net22 VPW n18 W=430.00n L=180.00n
MM9 net30 D net14 VPW n18 W=0.565u L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM23 net0152 cn net0157 VPW n18 W=430.00n L=180.00n
MM22 net0157 net0153 VSS VPW n18 W=430.00n L=180.00n
MM19 net0153 net0152 VSS VPW n18 W=430.00n L=180.00n
MM17 net0137 c net0152 VPW n18 W=430.00n L=180.00n
MM15 net0145 net0137 VSS VPW n18 W=430.00n L=180.00n
MM14 net18 c net0145 VPW n18 W=430.00n L=180.00n
MM11 net0137 net18 VSS VPW n18 W=430.00n L=180.00n
MM25 QN net0152 VSS VPW n18 W=560.00n L=180.00n
MM35 net94 RN net97 VNW p18 W=800.00n L=180.00n
MM24 QN net0152 VDD VNW p18 W=790.0n L=180.00n
MM21 net0224 net0153 VDD VNW p18 W=580.0n L=180.00n
MM20 net0152 c net0224 VNW p18 W=580.0n L=180.00n
MM18 net0153 net0152 VDD VNW p18 W=580.0n L=180.00n
MM16 net0137 cn net0152 VNW p18 W=580.0n L=180.00n
MM13 net18 cn net0212 VNW p18 W=570.0n L=180.00n
MM12 net0212 net0137 VDD VNW p18 W=570.0n L=180.00n
MM7 net97 SE VDD VNW p18 W=0.795u L=180.00n
MM0 net93 SI VDD VNW p18 W=490.0n L=180.00n
MM1 net94 SEN net93 VNW p18 W=490.0n L=180.00n
MM2 net94 D net97 VNW p18 W=0.795u L=180.00n
MM3 net18 c net94 VNW p18 W=710.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM10 net0137 net18 VDD VNW p18 W=570.0n L=180.00n
.ENDS SDGRNQNUHDV0P7
****Sub-Circuit for SDGRNQNUHDV1, Mon Jun 26 14:40:26 CST 2017****
.SUBCKT SDGRNQNUHDV1 CK D QN RN SE SI VDD VSS VNW VPW
MM34 net0152 RN VSS VPW n18 W=0.565u L=180.00n
MM6 net0148 SEN net0152 VPW n18 W=0.565u L=180.00n
MM4 net134 cn net0132 VPW n18 W=430.00n L=180.00n
MM5 net0140 SI VSS VPW n18 W=430.00n L=180.00n
MM8 net0132 SE net0140 VPW n18 W=430.00n L=180.00n
MM9 net0132 D net0148 VPW n18 W=0.565u L=180.00n
MM11 net0161 net134 VSS VPW n18 W=430.00n L=180.00n
MM14 net134 c net0153 VPW n18 W=430.00n L=180.00n
MM15 net0153 net0161 VSS VPW n18 W=430.00n L=180.00n
MM17 net0161 c net0123 VPW n18 W=430.00n L=180.00n
MM19 net0145 net0123 VSS VPW n18 W=430.00n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM22 net0141 net0145 VSS VPW n18 W=430.00n L=180.00n
MM23 net0123 cn net0141 VPW n18 W=430.00n L=180.00n
MM25 QN net0123 VSS VPW n18 W=720.00n L=180.00n
MM35 net0208 RN net0211 VNW p18 W=800.00n L=180.00n
MM7 net0211 SE VDD VNW p18 W=0.795u L=180.00n
MM0 net0215 SI VDD VNW p18 W=490.0n L=180.00n
MM1 net0208 SEN net0215 VNW p18 W=490.0n L=180.00n
MM2 net0208 D net0211 VNW p18 W=0.795u L=180.00n
MM3 net134 c net0208 VNW p18 W=710.00n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM21 net0212 net0145 VDD VNW p18 W=580.0n L=180.00n
MM10 net0161 net134 VDD VNW p18 W=570.0n L=180.00n
MM12 net0224 net0161 VDD VNW p18 W=570.0n L=180.00n
MM13 net134 cn net0224 VNW p18 W=570.0n L=180.00n
MM16 net0161 cn net0123 VNW p18 W=580.0n L=180.00n
MM18 net0145 net0123 VDD VNW p18 W=580.0n L=180.00n
MM20 net0123 c net0212 VNW p18 W=580.0n L=180.00n
MM24 QN net0123 VDD VNW p18 W=1.01u L=180.00n
.ENDS SDGRNQNUHDV1
****Sub-Circuit for SDGRNQNUHDV2, Mon Jun 26 14:40:26 CST 2017****
.SUBCKT SDGRNQNUHDV2 CK D QN RN SE SI VDD VSS VNW VPW
MM11 net0161 net134 VSS VPW n18 W=630.00n L=180.00n
MM14 net134 c net0153 VPW n18 W=410.00n L=180.00n
MM15 net0153 net0161 VSS VPW n18 W=410.00n L=180.00n
MM5 net0144 SI VSS VPW n18 W=430.00n L=180.00n
MM4 net134 cn net0152 VPW n18 W=490.00n L=180.00n
MM6 net0136 SEN net0132 VPW n18 W=0.565u L=180.00n
MM34 net0132 RN VSS VPW n18 W=0.565u L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM19 net0145 net0123 VSS VPW n18 W=430.00n L=180.00n
MM22 net0141 net0145 VSS VPW n18 W=430.00n L=180.00n
MM23 net0123 cn net0141 VPW n18 W=430.00n L=180.00n
MM9 net0152 D net0136 VPW n18 W=0.565u L=180.00n
MM8 net0152 SE net0144 VPW n18 W=430.00n L=180.00n
MM17 net0161 c net0123 VPW n18 W=630.00n L=180.00n
MM25 QN net0123 VSS VPW n18 W=1.44u L=180.00n
MM3 net134 c net0220 VNW p18 W=0.715u L=180.00n
MM2 net0220 D net0223 VNW p18 W=0.795u L=180.00n
MM1 net0220 SEN net0219 VNW p18 W=490.0n L=180.00n
MM0 net0219 SI VDD VNW p18 W=490.0n L=180.00n
MM7 net0223 SE VDD VNW p18 W=0.795u L=180.00n
MM35 net0220 RN net0223 VNW p18 W=800.00n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM21 net0212 net0145 VDD VNW p18 W=580.0n L=180.00n
MM24 QN net0123 VDD VNW p18 W=2.02u L=180.00n
MM10 net0161 net134 VDD VNW p18 W=0.89u L=180.00n
MM12 net0224 net0161 VDD VNW p18 W=580.0n L=180.00n
MM13 net134 cn net0224 VNW p18 W=580.0n L=180.00n
MM16 net0161 cn net0123 VNW p18 W=840.0n L=180.00n
MM18 net0145 net0123 VDD VNW p18 W=580.0n L=180.00n
MM20 net0123 c net0212 VNW p18 W=580.0n L=180.00n
.ENDS SDGRNQNUHDV2
****Sub-Circuit for SDGRSNQNUHDV0P7, Mon Jun 26 14:40:26 CST 2017****
.SUBCKT SDGRSNQNUHDV0P7 CK D QN RN SE SI SN VDD VSS VNW VPW
MM36 net0141 snn net0144 VPW n18 W=430.00n L=180.00n
MM37 snn SN VSS VPW n18 W=360.00n L=180.00n
MM6 net0144 RN net0149 VPW n18 W=0.565u L=180.00n
MM34 net0149 sen VSS VPW n18 W=0.565u L=180.00n
MM14 net18 c net0158 VPW n18 W=430.00n L=180.00n
MM11 net0150 net18 VSS VPW n18 W=430.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM31 sen SE VSS VPW n18 W=360.00n L=180.00n
MM9 net0141 D net0144 VPW n18 W=0.565u L=180.00n
MM8 net0141 SE net0201 VPW n18 W=430.00n L=180.00n
MM5 net0201 SI VSS VPW n18 W=430.00n L=180.00n
MM4 net18 cn net0141 VPW n18 W=430.00n L=180.00n
MM23 net0165 cn net0170 VPW n18 W=430.00n L=180.00n
MM22 net0170 net0166 VSS VPW n18 W=430.00n L=180.00n
MM19 net0166 net0165 VSS VPW n18 W=430.00n L=180.00n
MM17 net0150 c net0165 VPW n18 W=430.00n L=180.00n
MM15 net0158 net0150 VSS VPW n18 W=430.00n L=180.00n
MM25 QN net0165 VSS VPW n18 W=560.00n L=180.00n
MM38 snn SN VDD VNW p18 W=490.00n L=180.00n
MM24 QN net0165 VDD VNW p18 W=790.0n L=180.00n
MM21 net0245 net0166 VDD VNW p18 W=580.0n L=180.00n
MM20 net0165 c net0245 VNW p18 W=580.0n L=180.00n
MM18 net0166 net0165 VDD VNW p18 W=580.0n L=180.00n
MM16 net0150 cn net0165 VNW p18 W=580.0n L=180.00n
MM2 net0217 D net0236 VNW p18 W=0.795u L=180.00n
MM12 net0233 net0150 VDD VNW p18 W=570.0n L=180.00n
MM10 net0150 net18 VDD VNW p18 W=570.0n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM30 sen SE VDD VNW p18 W=490.00n L=180.00n
MM1 net0217 sen net0268 VNW p18 W=490.0n L=180.00n
MM0 net0268 SI VDD VNW p18 W=490.0n L=180.00n
MM7 net0220 SE VDD VNW p18 W=0.795u L=180.00n
MM35 net0217 RN net0220 VNW p18 W=490.00n L=180.00n
MM3 net18 c net0217 VNW p18 W=570.00n L=180.00n
MM39 net0236 snn net0220 VNW p18 W=0.795u L=180.00n
MM13 net18 cn net0233 VNW p18 W=570.0n L=180.00n
.ENDS SDGRSNQNUHDV0P7
****Sub-Circuit for SDGRSNQNUHDV1, Mon Jun 26 14:40:26 CST 2017****
.SUBCKT SDGRSNQNUHDV1 CK D QN RN SE SI SN VDD VSS VNW VPW
MM37 snn SN VSS VPW n18 W=360.00n L=180.00n
MM11 net0174 net134 VSS VPW n18 W=430.00n L=180.00n
MM14 net134 c net0166 VPW n18 W=430.00n L=180.00n
MM15 net0166 net0174 VSS VPW n18 W=430.00n L=180.00n
MM17 net0174 c net0165 VPW n18 W=430.00n L=180.00n
MM5 net0141 SI VSS VPW n18 W=430.00n L=180.00n
MM4 net134 cn net0157 VPW n18 W=430.00n L=180.00n
MM19 net0158 net0165 VSS VPW n18 W=430.00n L=180.00n
MM9 net0157 D net0160 VPW n18 W=0.565u L=180.00n
MM6 net0160 RN net0149 VPW n18 W=0.565u L=180.00n
MM34 net0149 sen VSS VPW n18 W=0.565u L=180.00n
MM8 net0157 SE net0141 VPW n18 W=430.00n L=180.00n
MM31 sen SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM22 net0154 net0158 VSS VPW n18 W=430.00n L=180.00n
MM23 net0165 cn net0154 VPW n18 W=430.00n L=180.00n
MM36 net0157 snn net0160 VPW n18 W=430.00n L=180.00n
MM25 QN net0165 VSS VPW n18 W=720.00n L=180.00n
MM38 snn SN VDD VNW p18 W=490.00n L=180.00n
MM35 net0233 RN net0240 VNW p18 W=490.00n L=180.00n
MM39 net0236 snn net0240 VNW p18 W=0.795u L=180.00n
MM2 net0233 D net0236 VNW p18 W=0.795u L=180.00n
MM7 net0240 SE VDD VNW p18 W=0.795u L=180.00n
MM1 net0233 sen net0228 VNW p18 W=490.0n L=180.00n
MM30 sen SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM21 net0135 net0158 VDD VNW p18 W=580.0n L=180.00n
MM10 net0174 net134 VDD VNW p18 W=570.0n L=180.00n
MM12 net0245 net0174 VDD VNW p18 W=570.0n L=180.00n
MM13 net134 cn net0245 VNW p18 W=570.0n L=180.00n
MM16 net0174 cn net0165 VNW p18 W=580.0n L=180.00n
MM0 net0228 SI VDD VNW p18 W=490.0n L=180.00n
MM3 net134 c net0233 VNW p18 W=570.00n L=180.00n
MM18 net0158 net0165 VDD VNW p18 W=580.0n L=180.00n
MM20 net0165 c net0135 VNW p18 W=580.0n L=180.00n
MM24 QN net0165 VDD VNW p18 W=1.01u L=180.00n
.ENDS SDGRSNQNUHDV1
****Sub-Circuit for SDGRSNQNUHDV2, Mon Jun 26 14:40:26 CST 2017****
.SUBCKT SDGRSNQNUHDV2 CK D QN RN SE SI SN VDD VSS VNW VPW
MM37 snn SN VSS VPW n18 W=360.00n L=180.00n
MM11 net0334 net134 VSS VPW n18 W=625.00n L=180.00n
MM14 net134 c net0326 VPW n18 W=410.00n L=180.00n
MM5 net0141 SI VSS VPW n18 W=430.00n L=180.00n
MM4 net134 cn net0157 VPW n18 W=430.00n L=180.00n
MM9 net0157 D net0160 VPW n18 W=0.565u L=180.00n
MM6 net0160 RN net0149 VPW n18 W=0.565u L=180.00n
MM34 net0149 sen VSS VPW n18 W=0.565u L=180.00n
MM8 net0157 SE net0141 VPW n18 W=430.00n L=180.00n
MM31 sen SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM17 net0334 c net0325 VPW n18 W=550.00n L=180.00n
MM19 net0318 net0325 VSS VPW n18 W=430.00n L=180.00n
MM22 net0314 net0318 VSS VPW n18 W=430.00n L=180.00n
MM23 net0325 cn net0314 VPW n18 W=430.00n L=180.00n
MM36 net0157 snn net0160 VPW n18 W=430.00n L=180.00n
MM15 net0326 net0334 VSS VPW n18 W=410.00n L=180.00n
MM25 QN net0325 VSS VPW n18 W=1.44u L=180.00n
MM38 snn SN VDD VNW p18 W=490.00n L=180.00n
MM35 net0233 RN net0240 VNW p18 W=490.00n L=180.00n
MM39 net0236 snn net0240 VNW p18 W=0.795u L=180.00n
MM2 net0233 D net0236 VNW p18 W=0.795u L=180.00n
MM7 net0240 SE VDD VNW p18 W=0.795u L=180.00n
MM1 net0233 sen net0228 VNW p18 W=490.0n L=180.00n
MM30 sen SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM18 net0318 net0325 VDD VNW p18 W=580.0n L=180.00n
MM20 net0325 c net0393 VNW p18 W=580.0n L=180.00n
MM21 net0393 net0318 VDD VNW p18 W=580.0n L=180.00n
MM24 QN net0325 VDD VNW p18 W=2.02u L=180.00n
MM10 net0334 net134 VDD VNW p18 W=860.00n L=180.00n
MM12 net0405 net0334 VDD VNW p18 W=580.0n L=180.00n
MM0 net0228 SI VDD VNW p18 W=490.0n L=180.00n
MM3 net134 c net0233 VNW p18 W=570.00n L=180.00n
MM13 net134 cn net0405 VNW p18 W=580.0n L=180.00n
MM16 net0334 cn net0325 VNW p18 W=800.00n L=180.00n
.ENDS SDGRSNQNUHDV2
.SUBCKT SDQNUHDV0P7 CK D QN SE SI VDD VSS VNW VPW
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM24 QN net101 VDD VNW p18 W=790.0n L=180.00n
MM21 net29 net94 VDD VNW p18 W=580.0n L=180.00n
MM20 net101 c net29 VNW p18 W=580.0n L=180.00n
MM18 net94 net101 VDD VNW p18 W=580.0n L=180.00n
MM16 net110 cn net101 VNW p18 W=580.0n L=180.00n
MM13 net130 cn net41 VNW p18 W=570.0n L=180.00n
MM12 net41 net110 VDD VNW p18 W=570.0n L=180.00n
MM10 net110 net130 VDD VNW p18 W=570.0n L=180.00n
MM3 net130 c net50 VNW p18 W=570.0n L=180.00n
MM2 net50 D net53 VNW p18 W=580.0n L=180.00n
MM1 net50 SEN net65 VNW p18 W=580.0n L=180.00n
MM0 net65 SI VDD VNW p18 W=580.0n L=180.00n
MM7 net53 SE VDD VNW p18 W=580.0n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM25 QN net101 VSS VPW n18 W=560.00n L=180.00n
MM23 net101 cn net90 VPW n18 W=430.00n L=180.00n
MM22 net90 net94 VSS VPW n18 W=430.00n L=180.00n
MM19 net94 net101 VSS VPW n18 W=430.00n L=180.00n
MM17 net110 c net101 VPW n18 W=430.00n L=180.00n
MM15 net102 net110 VSS VPW n18 W=430.00n L=180.00n
MM14 net130 c net102 VPW n18 W=430.00n L=180.00n
MM11 net110 net130 VSS VPW n18 W=430.00n L=180.00n
MM9 net114 D net118 VPW n18 W=430.00n L=180.00n
MM8 net114 SE net126 VPW n18 W=430.00n L=180.00n
MM5 net126 SI VSS VPW n18 W=430.00n L=180.00n
MM4 net130 cn net114 VPW n18 W=430.00n L=180.00n
MM6 net118 SEN VSS VPW n18 W=430.00n L=180.00n
.ENDS SDQNUHDV0P7
.SUBCKT SDQNUHDV1 CK D QN SE SI VDD VSS VNW VPW
MM6 net6 SEN VSS VPW n18 W=430.00n L=180.00n
MM4 net10 cn net22 VPW n18 W=430.00n L=180.00n
MM5 net14 SI VSS VPW n18 W=430.00n L=180.00n
MM8 net22 SE net14 VPW n18 W=430.00n L=180.00n
MM9 net22 D net6 VPW n18 W=430.00n L=180.00n
MM11 net26 net10 VSS VPW n18 W=430.00n L=180.00n
MM14 net10 c net34 VPW n18 W=430.00n L=180.00n
MM15 net34 net26 VSS VPW n18 W=430.00n L=180.00n
MM17 net26 c net41 VPW n18 W=430.00n L=180.00n
MM19 net42 net41 VSS VPW n18 W=430.00n L=180.00n
MM22 net46 net42 VSS VPW n18 W=430.00n L=180.00n
MM23 net41 cn net46 VPW n18 W=430.00n L=180.00n
MM25 QN net41 VSS VPW n18 W=720.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM7 net85 SE VDD VNW p18 W=580.0n L=180.00n
MM0 net81 SI VDD VNW p18 W=580.0n L=180.00n
MM1 net82 SEN net81 VNW p18 W=580.0n L=180.00n
MM2 net82 D net85 VNW p18 W=580.0n L=180.00n
MM3 net10 c net82 VNW p18 W=570.0n L=180.00n
MM10 net26 net10 VDD VNW p18 W=570.0n L=180.00n
MM12 net101 net26 VDD VNW p18 W=570.0n L=180.00n
MM13 net10 cn net101 VNW p18 W=570.0n L=180.00n
MM16 net26 cn net41 VNW p18 W=580.0n L=180.00n
MM18 net42 net41 VDD VNW p18 W=580.0n L=180.00n
MM20 net41 c net113 VNW p18 W=580.0n L=180.00n
MM21 net113 net42 VDD VNW p18 W=580.0n L=180.00n
MM24 QN net41 VDD VNW p18 W=1.01u L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
.ENDS SDQNUHDV1
.SUBCKT SDQNUHDV2 CK D QN SE SI VDD VSS VNW VPW
MM6 net6 SEN VSS VPW n18 W=560.00n L=180.00n
MM4 net10 cn net22 VPW n18 W=0.49u L=180.00n
MM5 net14 SI VSS VPW n18 W=560.00n L=180.00n
MM8 net22 SE net14 VPW n18 W=560.00n L=180.00n
MM9 net22 D net6 VPW n18 W=560.00n L=180.00n
MM11 net26 net10 VSS VPW n18 W=630.00n L=180.00n
MM14 net10 c net34 VPW n18 W=410.00n L=180.00n
MM15 net34 net26 VSS VPW n18 W=410.00n L=180.00n
MM17 net26 c net41 VPW n18 W=630.00n L=180.00n
MM19 net42 net41 VSS VPW n18 W=430.00n L=180.00n
MM22 net46 net42 VSS VPW n18 W=430.00n L=180.00n
MM23 net41 cn net46 VPW n18 W=430.00n L=180.00n
MM25 QN net41 VSS VPW n18 W=1.44u L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM7 net85 SE VDD VNW p18 W=790.0n L=180.00n
MM0 net81 SI VDD VNW p18 W=790.0n L=180.00n
MM1 net82 SEN net81 VNW p18 W=790.0n L=180.00n
MM2 net82 D net85 VNW p18 W=790.0n L=180.00n
MM3 net10 c net82 VNW p18 W=0.715u L=180.00n
MM10 net26 net10 VDD VNW p18 W=0.89u L=180.00n
MM12 net101 net26 VDD VNW p18 W=580.0n L=180.00n
MM13 net10 cn net101 VNW p18 W=580.0n L=180.00n
MM16 net26 cn net41 VNW p18 W=840.0n L=180.00n
MM18 net42 net41 VDD VNW p18 W=580.0n L=180.00n
MM20 net41 c net113 VNW p18 W=580.0n L=180.00n
MM21 net113 net42 VDD VNW p18 W=580.0n L=180.00n
MM24 QN net41 VDD VNW p18 W=2.02u L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
.ENDS SDQNUHDV2
.SUBCKT SDQUHDV0P7 CK D Q SE SI VDD VSS VNW VPW
MM6 net14 SEN VSS VPW n18 W=0.565u L=180.00n
MM4 net18 cn net30 VPW n18 W=0.575u L=180.00n
MM5 net22 SI VSS VPW n18 W=0.565u L=180.00n
MM8 net30 SE net22 VPW n18 W=0.565u L=180.00n
MM9 net30 D net14 VPW n18 W=0.565u L=180.00n
MM11 net34 net18 VSS VPW n18 W=0.56u L=180.00n
MM14 net18 c net42 VPW n18 W=0.405u L=180.00n
MM15 net42 net34 VSS VPW n18 W=0.405u L=180.00n
MM17 net6 net34 VSS VPW n18 W=0.635u L=180.00n
MM19 net46 net10 VSS VPW n18 W=0.435u L=180.00n
MM22 net50 net46 VSS VPW n18 W=0.435u L=180.00n
MM23 net10 cn net50 VPW n18 W=0.435u L=180.00n
MM25 Q net10 VSS VPW n18 W=0.57u L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM16 net10 c net6 VPW n18 W=0.635u L=180.00n
MM7 net97 SE VDD VNW p18 W=0.795u L=180.00n
MM0 net93 SI VDD VNW p18 W=0.8u L=180.00n
MM1 net94 SEN net93 VNW p18 W=0.8u L=180.00n
MM2 net94 D net97 VNW p18 W=0.795u L=180.00n
MM3 net18 c net94 VNW p18 W=0.715u L=180.00n
MM10 net34 net18 VDD VNW p18 W=0.69u L=180.00n
MM12 net113 net34 VDD VNW p18 W=0.59u L=180.00n
MM13 net18 cn net113 VNW p18 W=0.59u L=180.00n
MM32 net77 net34 VDD VNW p18 W=0.965u L=180.00n
MM18 net46 net10 VDD VNW p18 W=0.59u L=180.00n
MM20 net10 c net121 VNW p18 W=0.595u L=180.00n
MM21 net121 net46 VDD VNW p18 W=0.595u L=180.00n
MM24 Q net10 VDD VNW p18 W=0.8u L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM33 net10 cn net77 VNW p18 W=0.965u L=180.00n
.ENDS SDQUHDV0P7
.SUBCKT SDQUHDV1 CK D Q SE SI VDD VSS VNW VPW
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM24 Q net74 VDD VNW p18 W=1.01u L=180.00n
MM21 net37 net106 VDD VNW p18 W=0.595u L=180.00n
MM20 net74 c net37 VNW p18 W=0.595u L=180.00n
MM18 net106 net74 VDD VNW p18 W=0.59u L=180.00n
MM13 net134 cn net45 VNW p18 W=0.59u L=180.00n
MM12 net45 net118 VDD VNW p18 W=0.59u L=180.00n
MM10 net118 net134 VDD VNW p18 W=0.69u L=180.00n
MM3 net134 c net58 VNW p18 W=0.715u L=180.00n
MM2 net58 D net61 VNW p18 W=0.795u L=180.00n
MM1 net58 SEN net65 VNW p18 W=0.8u L=180.00n
MM0 net65 SI VDD VNW p18 W=0.8u L=180.00n
MM7 net61 SE VDD VNW p18 W=0.795u L=180.00n
MM16 net74 cn net13 VNW p18 W=0.965u L=180.00n
MM17 net13 net118 VDD VNW p18 W=0.965u L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM25 Q net74 VSS VPW n18 W=720.00n L=180.00n
MM23 net74 cn net102 VPW n18 W=0.435u L=180.00n
MM22 net102 net106 VSS VPW n18 W=0.435u L=180.00n
MM19 net106 net74 VSS VPW n18 W=0.435u L=180.00n
MM15 net110 net118 VSS VPW n18 W=0.405u L=180.00n
MM14 net134 c net110 VPW n18 W=0.405u L=180.00n
MM11 net118 net134 VSS VPW n18 W=0.56u L=180.00n
MM9 net122 D net138 VPW n18 W=0.565u L=180.00n
MM8 net122 SE net130 VPW n18 W=0.565u L=180.00n
MM5 net130 SI VSS VPW n18 W=0.565u L=180.00n
MM4 net134 cn net122 VPW n18 W=0.575u L=180.00n
MM6 net138 SEN VSS VPW n18 W=0.565u L=180.00n
MM32 net78 net118 VSS VPW n18 W=0.635u L=180.00n
MM33 net74 c net78 VPW n18 W=0.635u L=180.00n
.ENDS SDQUHDV1
.SUBCKT SDQUHDV2 CK D Q SE SI VDD VSS VNW VPW
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM24 Q net74 VDD VNW p18 W=2.02u L=180.00n
MM21 net37 net106 VDD VNW p18 W=0.595u L=180.00n
MM20 net74 c net37 VNW p18 W=0.595u L=180.00n
MM18 net106 net74 VDD VNW p18 W=0.59u L=180.00n
MM13 net134 cn net45 VNW p18 W=0.59u L=180.00n
MM12 net45 net118 VDD VNW p18 W=0.59u L=180.00n
MM10 net118 net134 VDD VNW p18 W=0.69u L=180.00n
MM3 net134 c net58 VNW p18 W=0.715u L=180.00n
MM2 net58 D net61 VNW p18 W=0.795u L=180.00n
MM1 net58 SEN net65 VNW p18 W=0.8u L=180.00n
MM0 net65 SI VDD VNW p18 W=0.8u L=180.00n
MM7 net61 SE VDD VNW p18 W=0.795u L=180.00n
MM16 net74 cn net13 VNW p18 W=0.965u L=180.00n
MM17 net13 net118 VDD VNW p18 W=0.965u L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM25 Q net74 VSS VPW n18 W=1.44u L=180.00n
MM23 net74 cn net102 VPW n18 W=0.435u L=180.00n
MM22 net102 net106 VSS VPW n18 W=0.435u L=180.00n
MM19 net106 net74 VSS VPW n18 W=0.435u L=180.00n
MM15 net110 net118 VSS VPW n18 W=0.405u L=180.00n
MM14 net134 c net110 VPW n18 W=0.405u L=180.00n
MM11 net118 net134 VSS VPW n18 W=560.00n L=180.00n
MM9 net122 D net138 VPW n18 W=0.565u L=180.00n
MM8 net122 SE net130 VPW n18 W=0.565u L=180.00n
MM5 net130 SI VSS VPW n18 W=0.565u L=180.00n
MM4 net134 cn net122 VPW n18 W=0.575u L=180.00n
MM6 net138 SEN VSS VPW n18 W=0.565u L=180.00n
MM32 net78 net118 VSS VPW n18 W=0.635u L=180.00n
MM33 net74 c net78 VPW n18 W=0.635u L=180.00n
.ENDS SDQUHDV2
.SUBCKT SDQUHDV3 CK D Q SE SI VDD VSS VNW VPW
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 c cn VDD VNW p18 W=420.00n L=180.00n
MM26 cn CK VDD VNW p18 W=250.00n L=180.00n
MM24 Q net74 VDD VNW p18 W=3.03u L=180.00n
MM21 net37 net106 VDD VNW p18 W=0.595u L=180.00n
MM20 net74 c net37 VNW p18 W=0.595u L=180.00n
MM18 net106 net74 VDD VNW p18 W=0.59u L=180.00n
MM13 net134 cn net45 VNW p18 W=0.59u L=180.00n
MM12 net45 net118 VDD VNW p18 W=0.59u L=180.00n
MM10 net118 net134 VDD VNW p18 W=0.69u L=180.00n
MM3 net134 c net58 VNW p18 W=0.715u L=180.00n
MM2 net58 D net61 VNW p18 W=0.795u L=180.00n
MM1 net58 SEN net65 VNW p18 W=0.8u L=180.00n
MM0 net65 SI VDD VNW p18 W=0.8u L=180.00n
MM7 net61 SE VDD VNW p18 W=0.795u L=180.00n
MM16 net74 cn net13 VNW p18 W=0.965u L=180.00n
MM17 net13 net118 VDD VNW p18 W=0.965u L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 c cn VSS VPW n18 W=250.00n L=180.00n
MM27 cn CK VSS VPW n18 W=420.00n L=180.00n
MM25 Q net74 VSS VPW n18 W=2.16u L=180.00n
MM23 net74 cn net102 VPW n18 W=0.435u L=180.00n
MM22 net102 net106 VSS VPW n18 W=0.435u L=180.00n
MM19 net106 net74 VSS VPW n18 W=0.435u L=180.00n
MM15 net110 net118 VSS VPW n18 W=0.405u L=180.00n
MM14 net134 c net110 VPW n18 W=0.405u L=180.00n
MM11 net118 net134 VSS VPW n18 W=560.00n L=180.00n
MM9 net122 D net138 VPW n18 W=0.565u L=180.00n
MM8 net122 SE net130 VPW n18 W=0.565u L=180.00n
MM5 net130 SI VSS VPW n18 W=0.565u L=180.00n
MM4 net134 cn net122 VPW n18 W=0.575u L=180.00n
MM6 net138 SEN VSS VPW n18 W=0.565u L=180.00n
MM32 net78 net118 VSS VPW n18 W=0.635u L=180.00n
MM33 net74 c net78 VPW n18 W=0.635u L=180.00n
.ENDS SDQUHDV3
.SUBCKT SDRNQUHDV0P7 CK D Q RDN SE SI VDD VSS VNW VPW
MM20 net7 RDN net_034 VPW n18 W=400.00n L=180.00n
MM21 net_034 net10 VSS VPW n18 W=400.00n L=180.00n
MM36 net_042 SEN VSS VPW n18 W=430.00n L=180.00n
MM35 net5 D net_042 VPW n18 W=430.00n L=180.00n
MM34 net_050 SI VSS VPW n18 W=430.00n L=180.00n
MM33 net5 SE net_050 VPW n18 W=430.00n L=180.00n
MM19 net9 cn net_074 VPW n18 W=0.42u L=180.00n
MM18 net_074 net4 VSS VPW n18 W=0.42u L=180.00n
MM14 net10 net6 VSS VPW n18 W=0.42u L=180.00n
MM12 net10 c net9 VPW n18 W=0.42u L=180.00n
MM10 Q net4 VSS VPW n18 W=560.00n L=180.00n
MM9 net4 net9 net_066 VPW n18 W=0.42u L=180.00n
MM8 net_066 RDN VSS VPW n18 W=0.42u L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM38 net7 c net6 VPW n18 W=790.00n L=180.00n
MM37 net5 cn net6 VPW n18 W=430.00n L=180.00n
MM23 net7 net10 VDD VNW p18 W=490.0n L=180.00n
MM22 net7 RDN VDD VNW p18 W=490.0n L=180.00n
MM32 net5 D net_0117 VNW p18 W=490.0n L=180.00n
MM31 net_0117 SE VDD VNW p18 W=490.0n L=180.00n
MM26 net_0129 SI VDD VNW p18 W=490.0n L=180.00n
MM25 net5 SEN net_0129 VNW p18 W=490.0n L=180.00n
MM17 net9 c net_0157 VNW p18 W=790.0n L=180.00n
MM16 net_0157 net4 VDD VNW p18 W=580.0n L=180.00n
MM15 net10 net6 VDD VNW p18 W=0.455u L=180.00n
MM13 net10 cn net9 VNW p18 W=0.825u L=180.00n
MM11 Q net4 VDD VNW p18 W=790.0n L=180.00n
MM3 net4 RDN VDD VNW p18 W=1060.0n L=180.00n
MM2 net4 net9 VDD VNW p18 W=1.01u L=180.00n
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM39 net7 cn net6 VNW p18 W=490.00n L=180.00n
MM40 net5 c net6 VNW p18 W=0.495u L=180.00n
.ENDS SDRNQUHDV0P7
.SUBCKT SDRNQUHDV1 CK D Q RDN SE SI VDD VSS VNW VPW
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM17 net9 c net_194 VNW p18 W=810.0n L=180.00n
MM16 net_194 net4 VDD VNW p18 W=580.0n L=180.00n
MM13 net10 cn net9 VNW p18 W=0.825u L=180.00n
MM11 Q net4 VDD VNW p18 W=1.01u L=180.00n
MM3 net4 RDN VDD VNW p18 W=1060.0n L=180.00n
MM2 net4 net9 VDD VNW p18 W=1.01u L=180.00n
MM39 net7 cn net6 VNW p18 W=490.00n L=180.00n
MM23 net7 net10 VDD VNW p18 W=490.0n L=180.00n
MM22 net7 RDN VDD VNW p18 W=490.0n L=180.00n
MM40 net5 c net6 VNW p18 W=0.495u L=180.00n
MM32 net5 D net_154 VNW p18 W=490.0n L=180.00n
MM31 net_154 SE VDD VNW p18 W=490.0n L=180.00n
MM26 net_142 SI VDD VNW p18 W=490.0n L=180.00n
MM25 net5 SEN net_142 VNW p18 W=490.0n L=180.00n
MM15 net10 net6 VDD VNW p18 W=0.455u L=180.00n
MM12 net10 c net9 VPW n18 W=0.42u L=180.00n
MM10 Q net4 VSS VPW n18 W=720.00n L=180.00n
MM9 net4 net9 net_243 VPW n18 W=0.42u L=180.00n
MM8 net_243 RDN VSS VPW n18 W=0.42u L=180.00n
MM38 net7 c net6 VPW n18 W=790.00n L=180.00n
MM20 net7 RDN net_231 VPW n18 W=400.00n L=180.00n
MM21 net_231 net10 VSS VPW n18 W=400.00n L=180.00n
MM37 net5 cn net6 VPW n18 W=430.00n L=180.00n
MM36 net_223 SEN VSS VPW n18 W=430.00n L=180.00n
MM35 net5 D net_223 VPW n18 W=430.00n L=180.00n
MM34 net_215 SI VSS VPW n18 W=430.00n L=180.00n
MM33 net5 SE net_215 VPW n18 W=430.00n L=180.00n
MM14 net10 net6 VSS VPW n18 W=0.42u L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM19 net9 cn net_259 VPW n18 W=0.42u L=180.00n
MM18 net_259 net4 VSS VPW n18 W=0.42u L=180.00n
.ENDS SDRNQUHDV1
.SUBCKT SDRNQUHDV2 CK D Q RDN SE SI VDD VSS VNW VPW
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM17 net9 c net_194 VNW p18 W=830.0n L=180.00n
MM16 net_194 net4 VDD VNW p18 W=580.0n L=180.00n
MM13 net10 cn net9 VNW p18 W=0.825u L=180.00n
MM11 Q net4 VDD VNW p18 W=2.02u L=180.00n
MM3 net4 RDN VDD VNW p18 W=1060.0n L=180.00n
MM2 net4 net9 VDD VNW p18 W=1.01u L=180.00n
MM39 net7 cn net6 VNW p18 W=490.00n L=180.00n
MM23 net7 net10 VDD VNW p18 W=490.0n L=180.00n
MM22 net7 RDN VDD VNW p18 W=490.0n L=180.00n
MM40 net5 c net6 VNW p18 W=0.495u L=180.00n
MM32 net5 D net_154 VNW p18 W=490.0n L=180.00n
MM31 net_154 SE VDD VNW p18 W=490.0n L=180.00n
MM26 net_142 SI VDD VNW p18 W=490.0n L=180.00n
MM25 net5 SEN net_142 VNW p18 W=490.0n L=180.00n
MM15 net10 net6 VDD VNW p18 W=0.455u L=180.00n
MM18 net_259 net4 VSS VPW n18 W=0.42u L=180.00n
MM12 net10 c net9 VPW n18 W=0.42u L=180.00n
MM10 Q net4 VSS VPW n18 W=1.44u L=180.00n
MM9 net4 net9 net_243 VPW n18 W=0.42u L=180.00n
MM8 net_243 RDN VSS VPW n18 W=0.42u L=180.00n
MM38 net7 c net6 VPW n18 W=790.00n L=180.00n
MM20 net7 RDN net_231 VPW n18 W=400.00n L=180.00n
MM21 net_231 net10 VSS VPW n18 W=400.00n L=180.00n
MM37 net5 cn net6 VPW n18 W=430.00n L=180.00n
MM36 net_223 SEN VSS VPW n18 W=430.00n L=180.00n
MM35 net5 D net_223 VPW n18 W=430.00n L=180.00n
MM34 net_215 SI VSS VPW n18 W=430.00n L=180.00n
MM33 net5 SE net_215 VPW n18 W=430.00n L=180.00n
MM14 net10 net6 VSS VPW n18 W=0.42u L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM19 net9 cn net_259 VPW n18 W=0.42u L=180.00n
.ENDS SDRNQUHDV2
.SUBCKT SDRNQUHDV3 CK D Q RDN SE SI VDD VSS VNW VPW
MM16 net_193 net4 VDD VNW p18 W=580.0n L=180.00n
MM13 net10 cn net9 VNW p18 W=825.000n L=180.00n
MM11 Q net4 VDD VNW p18 W=3.03u L=180.00n
MM3 net4 RDN VDD VNW p18 W=1.01u L=180.00n
MM2 net4 net9 VDD VNW p18 W=1.01u L=180.00n
MM39 net7 cn net6 VNW p18 W=495.00n L=180.00n
MM23 net7 net10 VDD VNW p18 W=490.0n L=180.00n
MM22 net7 RDN VDD VNW p18 W=495.00n L=180.00n
MM40 net5 c net6 VNW p18 W=0.495u L=180.00n
MM32 net5 D net_153 VNW p18 W=490.0n L=180.00n
MM31 net_153 SE VDD VNW p18 W=490.0n L=180.00n
MM26 net_141 SI VDD VNW p18 W=490.0n L=180.00n
MM25 net5 SEN net_141 VNW p18 W=490.0n L=180.00n
MM15 net10 net6 VDD VNW p18 W=0.455u L=180.00n
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM17 net9 c net_193 VNW p18 W=830.0n L=180.00n
MM8 net_258 RDN VSS VPW n18 W=0.42u L=180.00n
MM38 net7 c net6 VPW n18 W=790.00n L=180.00n
MM20 net7 RDN net_246 VPW n18 W=400.00n L=180.00n
MM21 net_246 net10 VSS VPW n18 W=400.00n L=180.00n
MM37 net5 cn net6 VPW n18 W=430.00n L=180.00n
MM36 net_238 SEN VSS VPW n18 W=430.00n L=180.00n
MM35 net5 D net_238 VPW n18 W=430.00n L=180.00n
MM34 net_230 SI VSS VPW n18 W=430.00n L=180.00n
MM33 net5 SE net_230 VPW n18 W=430.00n L=180.00n
MM14 net10 net6 VSS VPW n18 W=0.42u L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM18 net_274 net4 VSS VPW n18 W=0.42u L=180.00n
MM12 net10 c net9 VPW n18 W=0.42u L=180.00n
MM10 Q net4 VSS VPW n18 W=2.16u L=180.00n
MM9 net4 net9 net_258 VPW n18 W=0.42u L=180.00n
MM19 net9 cn net_274 VPW n18 W=0.42u L=180.00n
.ENDS SDRNQUHDV3
****Sub-Circuit for SDRQUHDV0P7, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT SDRQUHDV0P7 CK D Q RD SE SI VDD VSS VNW VPW
MM34 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM0 net075 D net091 VPW n18 W=0.565u L=180.00n
MM2 net083 SI VSS VPW n18 W=420.00n L=180.00n
MM1 net075 SE net083 VPW n18 W=420.00n L=180.00n
MM28 net091 SEN VSS VPW n18 W=0.565u L=180.00n
MM3 net17 cn net075 VPW n18 W=0.575u L=180.00n
MM22 Q net47 VSS VPW n18 W=560.00n L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=420.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM35 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM23 Q net47 VDD VNW p18 W=790.00n L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=790.00n L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
MM33 net0154 SE VDD VNW p18 W=0.795u L=180.00n
MM32 net0158 SI VDD VNW p18 W=420.0n L=180.00n
MM31 net0151 SEN net0158 VNW p18 W=420.0n L=180.00n
MM30 net0151 D net0154 VNW p18 W=0.795u L=180.00n
MM29 net17 c net0151 VNW p18 W=0.715u L=180.00n
.ENDS SDRQUHDV0P7
****Sub-Circuit for SDRQUHDV1, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT SDRQUHDV1 CK D Q RD SE SI VDD VSS VNW VPW
MM34 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM2 net083 SI VSS VPW n18 W=420.00n L=180.00n
MM1 net075 SE net083 VPW n18 W=420.00n L=180.00n
MM0 net075 D net091 VPW n18 W=0.565u L=180.00n
MM22 Q net47 VSS VPW n18 W=720.00n L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM28 net091 SEN VSS VPW n18 W=0.565u L=180.00n
MM3 net17 cn net075 VPW n18 W=0.575u L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=560.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM35 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM23 Q net47 VDD VNW p18 W=1.01u L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=1.01u L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
MM33 net0154 SE VDD VNW p18 W=0.795u L=180.00n
MM32 net0158 SI VDD VNW p18 W=420.0n L=180.00n
MM31 net0151 SEN net0158 VNW p18 W=420.0n L=180.00n
MM30 net0151 D net0154 VNW p18 W=0.795u L=180.00n
MM29 net17 c net0151 VNW p18 W=0.715u L=180.00n
.ENDS SDRQUHDV1
****Sub-Circuit for SDRQUHDV2, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT SDRQUHDV2 CK D Q RD SE SI VDD VSS VNW VPW
MM34 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM0 net075 D net091 VPW n18 W=0.565u L=180.00n
MM2 net083 SI VSS VPW n18 W=420.00n L=180.00n
MM1 net075 SE net083 VPW n18 W=420.00n L=180.00n
MM28 net091 SEN VSS VPW n18 W=0.565u L=180.00n
MM3 net17 cn net075 VPW n18 W=0.575u L=180.00n
MM22 Q net47 VSS VPW n18 W=1.44u L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=560.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM35 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM23 Q net47 VDD VNW p18 W=2.02u L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=1.01u L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
MM33 net0154 SE VDD VNW p18 W=0.795u L=180.00n
MM32 net0158 SI VDD VNW p18 W=420.0n L=180.00n
MM31 net0151 SEN net0158 VNW p18 W=420.0n L=180.00n
MM30 net0151 D net0154 VNW p18 W=0.795u L=180.00n
MM29 net17 c net0151 VNW p18 W=0.715u L=180.00n
.ENDS SDRQUHDV2
****Sub-Circuit for SDRQUHDV3, Tue Jun 13 08:55:59 CST 2017****
.SUBCKT SDRQUHDV3 CK D Q RD SE SI VDD VSS VNW VPW
MM34 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM22 Q net47 VSS VPW n18 W=2.16u L=180.00n
MM27 net44 RD VSS VPW n18 W=280.00n L=180.00n
MM17 net44 cn net45 VPW n18 W=280.00n L=180.00n
MM9 net53 net37 VSS VPW n18 W=280.00n L=180.00n
MM14 net37 c net44 VPW n18 W=300.00n L=180.00n
MM25 net37 RD VSS VPW n18 W=280.00n L=180.00n
MM6 net17 c net53 VPW n18 W=280.00n L=180.00n
MM18 net47 net44 VSS VPW n18 W=560.00n L=180.00n
MM4 net37 net17 VSS VPW n18 W=420.00n L=180.00n
MM16 net45 net47 VSS VPW n18 W=280.00n L=180.00n
MM12 c cn VSS VPW n18 W=280.00n L=180.00n
MM10 cn CK VSS VPW n18 W=420.00n L=180.00n
MM0 net091 D net075 VPW n18 W=0.565u L=180.00n
MM1 net091 SE net083 VPW n18 W=420.00n L=180.00n
MM2 net083 SI VSS VPW n18 W=420.00n L=180.00n
MM3 net17 cn net091 VPW n18 W=0.575u L=180.00n
MM28 net075 SEN VSS VPW n18 W=0.565u L=180.00n
MM35 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM23 Q net47 VDD VNW p18 W=3.03u L=180.00n
MM24 net80 RD VDD VNW p18 W=515.00n L=180.00n
MM21 net47 net44 VDD VNW p18 W=1.01u L=180.00n
MM26 net104 RD VDD VNW p18 W=280.00n L=180.00n
MM20 net44 c net100 VNW p18 W=280.00n L=180.00n
MM19 net100 net47 net104 VNW p18 W=280.00n L=180.00n
MM15 net37 cn net44 VNW p18 W=450.00n L=180.00n
MM8 net108 net37 VDD VNW p18 W=280.00n L=180.00n
MM7 net17 cn net108 VNW p18 W=280.00n L=180.00n
MM5 net37 net17 net80 VNW p18 W=515.00n L=180.00n
MM13 c cn VDD VNW p18 W=420.00n L=180.00n
MM11 cn CK VDD VNW p18 W=280.00n L=180.00n
MM29 net17 c net0159 VNW p18 W=0.715u L=180.00n
MM30 net0159 D net0162 VNW p18 W=0.795u L=180.00n
MM31 net0159 SEN net0158 VNW p18 W=420.0n L=180.00n
MM32 net0158 SI VDD VNW p18 W=420.0n L=180.00n
MM33 net0162 SE VDD VNW p18 W=0.795u L=180.00n
.ENDS SDRQUHDV3
.SUBCKT SDSNQUHDV0P7 CK D Q SDN SE SI VDD VSS VNW VPW
MM11 net_7 net_9 VDD VNW p18 W=0.765u L=180.00n
MM12 net_7 SDN VDD VNW p18 W=960.0n L=180.00n
MM43 net_7 c net_98 VNW p18 W=730.0n L=180.00n
MM44 net_117 cn net_98 VNW p18 W=0.74u L=180.00n
MM9 net_9 net_98 VDD VNW p18 W=0.95u L=180.00n
MM40 net_115 cn net6 VNW p18 W=495.00n L=180.00n
MM39 net7 c net6 VNW p18 W=0.495u L=180.00n
MM22 net_115 net_117 VDD VNW p18 W=0.495u L=180.00n
MM25 net7 SEN net_42 VNW p18 W=490.0n L=180.00n
MM26 net_42 SI VDD VNW p18 W=490.0n L=180.00n
MM31 net_54 SE VDD VNW p18 W=490.0n L=180.00n
MM32 net7 D net_54 VNW p18 W=490.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM3 Q net_9 VDD VNW p18 W=0.71u L=180.00n
MM15 net_117 net6 VDD VNW p18 W=0.495u L=180.00n
MM14 net_117 SDN VDD VNW p18 W=0.495u L=180.00n
MM10 net_79 net_9 VSS VPW n18 W=430.00n L=180.00n
MM13 net_7 SDN net_79 VPW n18 W=400.00n L=180.00n
MM20 net_117 net6 net_91 VPW n18 W=400.00n L=180.00n
MM21 net_91 SDN VSS VPW n18 W=400.00n L=180.00n
MM41 net_7 cn net_98 VPW n18 W=400.00n L=180.00n
MM42 net_117 c net_98 VPW n18 W=0.39u L=180.00n
MM8 net_9 net_98 VSS VPW n18 W=510.00n L=180.00n
MM37 net_115 c net6 VPW n18 W=0.385u L=180.00n
MM38 net7 cn net6 VPW n18 W=0.43u L=180.00n
MM29 net_115 net_117 VSS VPW n18 W=430.00n L=180.00n
MM33 net7 SE net_123 VPW n18 W=430.00n L=180.00n
MM34 net_123 SI VSS VPW n18 W=430.00n L=180.00n
MM35 net7 D net_131 VPW n18 W=430.00n L=180.00n
MM36 net_131 SEN VSS VPW n18 W=430.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM2 Q net_9 VSS VPW n18 W=560.00n L=180.00n
.ENDS SDSNQUHDV0P7
.SUBCKT SDSNQUHDV1 CK D Q SDN SE SI VDD VSS VNW VPW
MM10 net_211 net_183 VSS VPW n18 W=430.00n L=180.00n
MM13 net_203 SDN net_211 VPW n18 W=400.00n L=180.00n
MM41 net_203 cn net_182 VPW n18 W=400.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM2 Q net_183 VSS VPW n18 W=720.00n L=180.00n
MM8 net_183 net_182 VSS VPW n18 W=510.00n L=180.00n
MM42 net_167 c net_182 VPW n18 W=0.39u L=180.00n
MM37 net_175 c net6 VPW n18 W=0.385u L=180.00n
MM29 net_175 net_167 VSS VPW n18 W=430.00n L=180.00n
MM20 net_167 net6 net_163 VPW n18 W=400.00n L=180.00n
MM21 net_163 SDN VSS VPW n18 W=400.00n L=180.00n
MM33 net7 SE net_155 VPW n18 W=430.00n L=180.00n
MM34 net_155 SI VSS VPW n18 W=430.00n L=180.00n
MM35 net7 D net_147 VPW n18 W=430.00n L=180.00n
MM36 net_147 SEN VSS VPW n18 W=430.00n L=180.00n
MM38 net7 cn net6 VPW n18 W=0.43u L=180.00n
MM15 net_167 net6 VDD VNW p18 W=0.495u L=180.00n
MM14 net_167 SDN VDD VNW p18 W=0.495u L=180.00n
MM25 net7 SEN net_234 VNW p18 W=490.0n L=180.00n
MM26 net_234 SI VDD VNW p18 W=490.0n L=180.00n
MM31 net_222 SE VDD VNW p18 W=490.0n L=180.00n
MM32 net7 D net_222 VNW p18 W=490.0n L=180.00n
MM39 net7 c net6 VNW p18 W=0.495u L=180.00n
MM11 net_203 net_183 VDD VNW p18 W=0.765u L=180.00n
MM12 net_203 SDN VDD VNW p18 W=960.0n L=180.00n
MM43 net_203 c net_182 VNW p18 W=730.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM3 Q net_183 VDD VNW p18 W=1.01u L=180.00n
MM9 net_183 net_182 VDD VNW p18 W=0.95u L=180.00n
MM44 net_167 cn net_182 VNW p18 W=0.74u L=180.00n
MM40 net_175 cn net6 VNW p18 W=495.00n L=180.00n
MM22 net_175 net_167 VDD VNW p18 W=0.495u L=180.00n
.ENDS SDSNQUHDV1
.SUBCKT SDSNQUHDV2 CK D Q SDN SE SI VDD VSS VNW VPW
MM39 net7 c net6 VNW p18 W=0.495u L=180.00n
MM32 net7 D net_210 VNW p18 W=490.0n L=180.00n
MM31 net_210 SE VDD VNW p18 W=490.0n L=180.00n
MM26 net_198 SI VDD VNW p18 W=490.0n L=180.00n
MM25 net7 SEN net_198 VNW p18 W=490.0n L=180.00n
MM14 net_259 SDN VDD VNW p18 W=0.495u L=180.00n
MM15 net_259 net6 VDD VNW p18 W=0.495u L=180.00n
MM22 net_251 net_259 VDD VNW p18 W=0.495u L=180.00n
MM40 net_251 cn net6 VNW p18 W=495.00n L=180.00n
MM44 net_259 cn net_250 VNW p18 W=0.74u L=180.00n
MM9 net_243 net_250 VDD VNW p18 W=0.95u L=180.00n
MM3 Q net_243 VDD VNW p18 W=2.02u L=180.00n
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM43 net_223 c net_250 VNW p18 W=730.0n L=180.00n
MM12 net_223 SDN VDD VNW p18 W=960.0n L=180.00n
MM11 net_223 net_243 VDD VNW p18 W=0.765u L=180.00n
MM35 net7 D net_279 VPW n18 W=430.00n L=180.00n
MM34 net_271 SI VSS VPW n18 W=430.00n L=180.00n
MM33 net7 SE net_271 VPW n18 W=430.00n L=180.00n
MM21 net_263 SDN VSS VPW n18 W=400.00n L=180.00n
MM20 net_259 net6 net_263 VPW n18 W=400.00n L=180.00n
MM29 net_251 net_259 VSS VPW n18 W=430.00n L=180.00n
MM37 net_251 c net6 VPW n18 W=0.385u L=180.00n
MM42 net_259 c net_250 VPW n18 W=0.39u L=180.00n
MM8 net_243 net_250 VSS VPW n18 W=510.00n L=180.00n
MM2 Q net_243 VSS VPW n18 W=1.44u L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM41 net_223 cn net_250 VPW n18 W=400.00n L=180.00n
MM13 net_223 SDN net_215 VPW n18 W=400.00n L=180.00n
MM10 net_215 net_243 VSS VPW n18 W=430.00n L=180.00n
MM38 net7 cn net6 VPW n18 W=0.43u L=180.00n
MM36 net_279 SEN VSS VPW n18 W=430.00n L=180.00n
.ENDS SDSNQUHDV2
.SUBCKT SDSNQUHDV3 CK D Q SDN SE SI VDD VSS VNW VPW
MM31 net_208 SE VDD VNW p18 W=490.0n L=180.00n
MM26 net_196 SI VDD VNW p18 W=490.0n L=180.00n
MM25 net7 SEN net_196 VNW p18 W=490.0n L=180.00n
MM14 net_265 SDN VDD VNW p18 W=0.495u L=180.00n
MM15 net_265 net6 VDD VNW p18 W=0.495u L=180.00n
MM22 net_257 net_265 VDD VNW p18 W=0.495u L=180.00n
MM40 net_257 cn net6 VNW p18 W=495.00n L=180.00n
MM44 net_265 cn net_256 VNW p18 W=0.74u L=180.00n
MM9 net_249 net_256 VDD VNW p18 W=0.95u L=180.00n
MM3 Q net_249 VDD VNW p18 W=3.03u L=180.00n
MM1 c cn VDD VNW p18 W=420.00n L=180.00n
MM7 SEN SE VDD VNW p18 W=490.0n L=180.00n
MM5 cn CK VDD VNW p18 W=250.00n L=180.00n
MM43 net_229 c net_256 VNW p18 W=730.0n L=180.00n
MM12 net_229 SDN VDD VNW p18 W=960.0n L=180.00n
MM11 net_229 net_249 VDD VNW p18 W=0.765u L=180.00n
MM39 net7 c net6 VNW p18 W=0.495u L=180.00n
MM32 net7 D net_208 VNW p18 W=490.0n L=180.00n
MM36 net_213 SEN VSS VPW n18 W=430.00n L=180.00n
MM35 net7 D net_213 VPW n18 W=430.00n L=180.00n
MM34 net_277 SI VSS VPW n18 W=430.00n L=180.00n
MM33 net7 SE net_277 VPW n18 W=430.00n L=180.00n
MM21 net_269 SDN VSS VPW n18 W=400.00n L=180.00n
MM20 net_265 net6 net_269 VPW n18 W=400.00n L=180.00n
MM29 net_257 net_265 VSS VPW n18 W=430.00n L=180.00n
MM37 net_257 c net6 VPW n18 W=0.385u L=180.00n
MM42 net_265 c net_256 VPW n18 W=0.39u L=180.00n
MM8 net_249 net_256 VSS VPW n18 W=510.00n L=180.00n
MM2 Q net_249 VSS VPW n18 W=2.16u L=180.00n
MM0 c cn VSS VPW n18 W=250.00n L=180.00n
MM6 SEN SE VSS VPW n18 W=430.00n L=180.00n
MM4 cn CK VSS VPW n18 W=420.00n L=180.00n
MM41 net_229 cn net_256 VPW n18 W=400.00n L=180.00n
MM13 net_229 SDN net_221 VPW n18 W=400.00n L=180.00n
MM10 net_221 net_249 VSS VPW n18 W=430.00n L=180.00n
MM38 net7 cn net6 VPW n18 W=0.43u L=180.00n
.ENDS SDSNQUHDV3
.SUBCKT SDSRNQUHDV1 CK D Q RDN SDN SE SI VDD VSS VNW VPW
MM40 net0163 SEN net082 VNW p18 W=0.36u L=180.00n
MM29 net0163 D net61 VNW p18 W=0.69u L=180.00n
MM41 net082 SI VDD VNW p18 W=0.36u L=180.00n
MM46 SEN SE VDD VNW p18 W=0.485u L=180.00n
MM44 net0163 c net108 VNW p18 W=0.42u L=180.00n
MM30 net101 SDN VDD VNW p18 W=0.37u L=180.00n
MM32 net108 cn net88 VNW p18 W=0.42u L=180.00n
MM21 net88 net101 VDD VNW p18 W=0.42u L=180.00n
MM20 net88 RDN VDD VNW p18 W=0.42u L=180.00n
MM14 net101 cn net100 VNW p18 W=0.425u L=180.00n
MM10 net101 net108 VDD VNW p18 W=0.42u L=180.00n
MM6 c cn VDD VNW p18 W=420.00n L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM0 net61 SE VDD VNW p18 W=0.69u L=180.00n
MM16 net112 RDN VDD VNW p18 W=0.42u L=180.00n
MM17 net112 net100 VDD VNW p18 W=0.42u L=180.00n
MM5 Q net112 VDD VNW p18 W=1.01u L=180.00n
MM34 net0204 net112 VDD VNW p18 W=0.42u L=180.00n
MM35 net0204 SDN VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net0204 VNW p18 W=0.425u L=180.00n
MM43 net0155 SI VSS VPW n18 W=0.445u L=180.00n
MM42 net0163 SE net0155 VPW n18 W=0.445u L=180.00n
MM47 SEN SE VSS VPW n18 W=0.52u L=180.00n
MM37 net100 cn net0264 VPW n18 W=0.42u L=180.00n
MM38 net0264 SDN net0260 VPW n18 W=0.42u L=180.00n
MM33 net108 c net0292 VPW n18 W=0.445u L=180.00n
MM45 net0163 cn net108 VPW n18 W=0.445u L=180.00n
MM31 net0276 net108 VSS VPW n18 W=0.49u L=180.00n
MM28 net0163 D net0320 VPW n18 W=0.445u L=180.00n
MM39 net0260 net112 VSS VPW n18 W=0.42u L=180.00n
MM1 net0320 SEN VSS VPW n18 W=0.445u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM3 cn CK VSS VPW n18 W=420.00n L=180.00n
MM19 net112 net100 net77 VPW n18 W=0.53u L=180.00n
MM18 net77 RDN VSS VPW n18 W=0.53u L=180.00n
MM23 net0292 RDN net93 VPW n18 W=0.445u L=180.00n
MM22 net93 net101 VSS VPW n18 W=0.445u L=180.00n
MM15 net101 c net100 VPW n18 W=0.42u L=180.00n
MM12 net101 SDN net0276 VPW n18 W=0.49u L=180.00n
MM4 Q net112 VSS VPW n18 W=0.72u L=180.00n
.ENDS SDSRNQUHDV1
.SUBCKT SDSRNQUHDV2 CK D Q RDN SDN SE SI VDD VSS VNW VPW
MM40 net0163 SEN net082 VNW p18 W=0.36u L=180.00n
MM29 net0163 D net61 VNW p18 W=0.69u L=180.00n
MM41 net082 SI VDD VNW p18 W=0.36u L=180.00n
MM46 SEN SE VDD VNW p18 W=0.485u L=180.00n
MM44 net0163 c net108 VNW p18 W=0.42u L=180.00n
MM30 net101 SDN VDD VNW p18 W=0.37u L=180.00n
MM32 net108 cn net88 VNW p18 W=0.42u L=180.00n
MM21 net88 net101 VDD VNW p18 W=0.42u L=180.00n
MM20 net88 RDN VDD VNW p18 W=0.42u L=180.00n
MM14 net101 cn net100 VNW p18 W=0.425u L=180.00n
MM10 net101 net108 VDD VNW p18 W=0.42u L=180.00n
MM6 c cn VDD VNW p18 W=420.00n L=180.00n
MM2 cn CK VDD VNW p18 W=250.00n L=180.00n
MM0 net61 SE VDD VNW p18 W=0.69u L=180.00n
MM16 net112 RDN VDD VNW p18 W=0.42u L=180.00n
MM17 net112 net100 VDD VNW p18 W=0.42u L=180.00n
MM5 Q net112 VDD VNW p18 W=2.02u L=180.00n
MM34 net0204 net112 VDD VNW p18 W=0.42u L=180.00n
MM35 net0204 SDN VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net0204 VNW p18 W=0.425u L=180.00n
MM43 net0155 SI VSS VPW n18 W=0.445u L=180.00n
MM42 net0163 SE net0155 VPW n18 W=0.445u L=180.00n
MM47 SEN SE VSS VPW n18 W=0.52u L=180.00n
MM37 net100 cn net0264 VPW n18 W=0.42u L=180.00n
MM38 net0264 SDN net0260 VPW n18 W=0.42u L=180.00n
MM33 net108 c net0292 VPW n18 W=0.445u L=180.00n
MM45 net0163 cn net108 VPW n18 W=0.445u L=180.00n
MM31 net0276 net108 VSS VPW n18 W=0.49u L=180.00n
MM28 net0163 D net0320 VPW n18 W=0.445u L=180.00n
MM39 net0260 net112 VSS VPW n18 W=0.42u L=180.00n
MM1 net0320 SEN VSS VPW n18 W=0.445u L=180.00n
MM7 c cn VSS VPW n18 W=250.00n L=180.00n
MM3 cn CK VSS VPW n18 W=420.00n L=180.00n
MM19 net112 net100 net77 VPW n18 W=0.53u L=180.00n
MM18 net77 RDN VSS VPW n18 W=0.53u L=180.00n
MM23 net0292 RDN net93 VPW n18 W=0.445u L=180.00n
MM22 net93 net101 VSS VPW n18 W=0.445u L=180.00n
MM15 net101 c net100 VPW n18 W=0.42u L=180.00n
MM12 net101 SDN net0276 VPW n18 W=0.49u L=180.00n
MM4 Q net112 VSS VPW n18 W=1.44u L=180.00n
.ENDS SDSRNQUHDV2
.SUBCKT SNDQUHDV0P7 CKN D Q SE SI VDD VSS VNW VPW
MM33 net74 cn net9 VNW p18 W=580.0n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 cn c VDD VNW p18 W=250.00n L=180.00n
MM26 c CKN VDD VNW p18 W=420.00n L=180.00n
MM24 Q net74 VDD VNW p18 W=790.0n L=180.00n
MM21 net33 net102 VDD VNW p18 W=580.0n L=180.00n
MM20 net74 c net33 VNW p18 W=580.0n L=180.00n
MM18 net102 net74 VDD VNW p18 W=580.0n L=180.00n
MM32 net9 net118 VDD VNW p18 W=0.52u L=180.00n
MM13 net134 cn net45 VNW p18 W=0.52u L=180.00n
MM12 net45 net118 VDD VNW p18 W=0.52u L=180.00n
MM10 net118 net134 VDD VNW p18 W=0.52u L=180.00n
MM3 net134 c net58 VNW p18 W=570.0n L=180.00n
MM2 net58 D net61 VNW p18 W=580.0n L=180.00n
MM1 net58 SI net65 VNW p18 W=580.0n L=180.00n
MM0 net65 SEN VDD VNW p18 W=580.0n L=180.00n
MM7 net61 SE VDD VNW p18 W=580.0n L=180.00n
MM16 net74 c net106 VPW n18 W=430.00n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 cn c VSS VPW n18 W=420.00n L=180.00n
MM27 c CKN VSS VPW n18 W=250.00n L=180.00n
MM25 Q net74 VSS VPW n18 W=560.00n L=180.00n
MM23 net74 cn net98 VPW n18 W=430.00n L=180.00n
MM22 net98 net102 VSS VPW n18 W=430.00n L=180.00n
MM19 net102 net74 VSS VPW n18 W=430.00n L=180.00n
MM17 net106 net118 VSS VPW n18 W=430.00n L=180.00n
MM15 net110 net118 VSS VPW n18 W=430.00n L=180.00n
MM14 net134 c net110 VPW n18 W=430.00n L=180.00n
MM11 net118 net134 VSS VPW n18 W=430.00n L=180.00n
MM9 net122 D net138 VPW n18 W=430.00n L=180.00n
MM8 net122 SI net130 VPW n18 W=430.00n L=180.00n
MM5 net130 SE VSS VPW n18 W=430.00n L=180.00n
MM4 net134 cn net122 VPW n18 W=430.00n L=180.00n
MM6 net138 SEN VSS VPW n18 W=430.00n L=180.00n
.ENDS SNDQUHDV0P7
.SUBCKT SNDQUHDV1 CKN D Q SE SI VDD VSS VNW VPW
MM6 net6 SEN VSS VPW n18 W=430.00n L=180.00n
MM4 net10 cn net22 VPW n18 W=430.00n L=180.00n
MM5 net14 SE VSS VPW n18 W=430.00n L=180.00n
MM8 net22 SI net14 VPW n18 W=430.00n L=180.00n
MM9 net22 D net6 VPW n18 W=430.00n L=180.00n
MM11 net26 net10 VSS VPW n18 W=430.00n L=180.00n
MM14 net10 c net34 VPW n18 W=430.00n L=180.00n
MM15 net34 net26 VSS VPW n18 W=430.00n L=180.00n
MM17 net38 net26 VSS VPW n18 W=430.00n L=180.00n
MM19 net42 net70 VSS VPW n18 W=430.00n L=180.00n
MM22 net46 net42 VSS VPW n18 W=430.00n L=180.00n
MM23 net70 cn net46 VPW n18 W=430.00n L=180.00n
MM25 Q net70 VSS VPW n18 W=720.00n L=180.00n
MM27 c CKN VSS VPW n18 W=250.00n L=180.00n
MM29 cn c VSS VPW n18 W=420.00n L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM16 net70 c net38 VPW n18 W=430.00n L=180.00n
MM7 net89 SE VDD VNW p18 W=580.0n L=180.00n
MM0 net85 SEN VDD VNW p18 W=580.0n L=180.00n
MM1 net86 SI net85 VNW p18 W=580.0n L=180.00n
MM2 net86 D net89 VNW p18 W=580.0n L=180.00n
MM3 net10 c net86 VNW p18 W=570.0n L=180.00n
MM10 net26 net10 VDD VNW p18 W=0.52u L=180.00n
MM12 net105 net26 VDD VNW p18 W=0.52u L=180.00n
MM13 net10 cn net105 VNW p18 W=0.52u L=180.00n
MM32 net141 net26 VDD VNW p18 W=0.52u L=180.00n
MM18 net42 net70 VDD VNW p18 W=580.0n L=180.00n
MM20 net70 c net117 VNW p18 W=580.0n L=180.00n
MM21 net117 net42 VDD VNW p18 W=580.0n L=180.00n
MM24 Q net70 VDD VNW p18 W=1.01u L=180.00n
MM26 c CKN VDD VNW p18 W=420.00n L=180.00n
MM28 cn c VDD VNW p18 W=250.00n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM33 net70 cn net141 VNW p18 W=580.0n L=180.00n
.ENDS SNDQUHDV1
.SUBCKT SNDQUHDV2 CKN D Q SE SI VDD VSS VNW VPW
MM33 net74 cn net9 VNW p18 W=950.0n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 cn c VDD VNW p18 W=250.00n L=180.00n
MM26 c CKN VDD VNW p18 W=420.00n L=180.00n
MM24 Q net74 VDD VNW p18 W=2.02u L=180.00n
MM21 net33 net102 VDD VNW p18 W=580.0n L=180.00n
MM20 net74 c net33 VNW p18 W=580.0n L=180.00n
MM18 net102 net74 VDD VNW p18 W=580.0n L=180.00n
MM32 net9 net118 VDD VNW p18 W=950.0n L=180.00n
MM13 net134 cn net45 VNW p18 W=580.0n L=180.00n
MM12 net45 net118 VDD VNW p18 W=580.0n L=180.00n
MM10 net118 net134 VDD VNW p18 W=790.0n L=180.00n
MM3 net134 c net58 VNW p18 W=0.74u L=180.00n
MM2 net58 D net61 VNW p18 W=790.0n L=180.00n
MM1 net58 SI net65 VNW p18 W=790.0n L=180.00n
MM0 net65 SEN VDD VNW p18 W=0.58u L=180.00n
MM7 net61 SE VDD VNW p18 W=790.0n L=180.00n
MM16 net74 c net106 VPW n18 W=0.43u L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 cn c VSS VPW n18 W=420.00n L=180.00n
MM27 c CKN VSS VPW n18 W=250.00n L=180.00n
MM25 Q net74 VSS VPW n18 W=1.44u L=180.00n
MM23 net74 cn net98 VPW n18 W=430.00n L=180.00n
MM22 net98 net102 VSS VPW n18 W=430.00n L=180.00n
MM19 net102 net74 VSS VPW n18 W=430.00n L=180.00n
MM17 net106 net118 VSS VPW n18 W=0.43u L=180.00n
MM15 net110 net118 VSS VPW n18 W=410.00n L=180.00n
MM14 net134 c net110 VPW n18 W=0.36u L=180.00n
MM11 net118 net134 VSS VPW n18 W=560.00n L=180.00n
MM9 net122 D net138 VPW n18 W=560.00n L=180.00n
MM8 net122 SI net130 VPW n18 W=560.00n L=180.00n
MM5 net130 SE VSS VPW n18 W=0.515u L=180.00n
MM4 net134 cn net122 VPW n18 W=430.00n L=180.00n
MM6 net138 SEN VSS VPW n18 W=560.00n L=180.00n
.ENDS SNDQUHDV2
.SUBCKT SNDQUHDV3 CKN D Q SE SI VDD VSS VNW VPW
MM33 net263 cn net198 VNW p18 W=950.0n L=180.00n
MM30 SEN SE VDD VNW p18 W=0.95u L=180.00n
MM28 cn c VDD VNW p18 W=250.00n L=180.00n
MM26 c CKN VDD VNW p18 W=420.00n L=180.00n
MM24 Q net263 VDD VNW p18 W=3.03u L=180.00n
MM21 net174 net235 VDD VNW p18 W=580.0n L=180.00n
MM20 net263 c net174 VNW p18 W=580.0n L=180.00n
MM18 net235 net263 VDD VNW p18 W=580.0n L=180.00n
MM32 net198 net219 VDD VNW p18 W=950.0n L=180.00n
MM13 net203 cn net162 VNW p18 W=580.0n L=180.00n
MM12 net162 net219 VDD VNW p18 W=580.0n L=180.00n
MM10 net219 net203 VDD VNW p18 W=790.0n L=180.00n
MM3 net203 c net143 VNW p18 W=0.74u L=180.00n
MM2 net143 D net146 VNW p18 W=790.0n L=180.00n
MM1 net143 SI net142 VNW p18 W=790.0n L=180.00n
MM0 net142 SEN VDD VNW p18 W=0.58u L=180.00n
MM7 net146 SE VDD VNW p18 W=790.0n L=180.00n
MM22 net239 net235 VSS VPW n18 W=430.00n L=180.00n
MM19 net235 net263 VSS VPW n18 W=430.00n L=180.00n
MM17 net231 net219 VSS VPW n18 W=0.43u L=180.00n
MM15 net227 net219 VSS VPW n18 W=410.00n L=180.00n
MM14 net203 c net227 VPW n18 W=0.36u L=180.00n
MM11 net219 net203 VSS VPW n18 W=560.00n L=180.00n
MM9 net215 D net199 VPW n18 W=560.00n L=180.00n
MM8 net215 SI net207 VPW n18 W=560.00n L=180.00n
MM5 net207 SE VSS VPW n18 W=0.515u L=180.00n
MM4 net203 cn net215 VPW n18 W=430.00n L=180.00n
MM6 net199 SEN VSS VPW n18 W=560.00n L=180.00n
MM16 net263 c net231 VPW n18 W=0.43u L=180.00n
MM31 SEN SE VSS VPW n18 W=720.00n L=180.00n
MM29 cn c VSS VPW n18 W=420.00n L=180.00n
MM27 c CKN VSS VPW n18 W=250.00n L=180.00n
MM25 Q net263 VSS VPW n18 W=2.16u L=180.00n
MM23 net263 cn net239 VPW n18 W=430.00n L=180.00n
.ENDS SNDQUHDV3
.SUBCKT SNDSRNQUHDV1 CKN D Q RDN SDN SE SI VDD VSS VNW VPW
MM40 net0163 SEN net082 VNW p18 W=0.36u L=180.00n
MM29 net0163 D net61 VNW p18 W=0.69u L=180.00n
MM41 net082 SI VDD VNW p18 W=0.36u L=180.00n
MM46 SEN SE VDD VNW p18 W=0.485u L=180.00n
MM44 net0163 c net108 VNW p18 W=0.42u L=180.00n
MM30 net101 SDN VDD VNW p18 W=0.37u L=180.00n
MM32 net108 cn net88 VNW p18 W=0.42u L=180.00n
MM21 net88 net101 VDD VNW p18 W=0.42u L=180.00n
MM20 net88 RDN VDD VNW p18 W=0.42u L=180.00n
MM14 net101 cn net100 VNW p18 W=0.425u L=180.00n
MM10 net101 net108 VDD VNW p18 W=0.42u L=180.00n
MM6 cn c VDD VNW p18 W=250.00n L=180.00n
MM2 c CKN VDD VNW p18 W=420.00n L=180.00n
MM0 net61 SE VDD VNW p18 W=0.69u L=180.00n
MM16 net112 RDN VDD VNW p18 W=0.42u L=180.00n
MM17 net112 net100 VDD VNW p18 W=0.42u L=180.00n
MM5 Q net112 VDD VNW p18 W=1.01u L=180.00n
MM34 net0204 net112 VDD VNW p18 W=0.42u L=180.00n
MM35 net0204 SDN VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net0204 VNW p18 W=0.425u L=180.00n
MM43 net0155 SI VSS VPW n18 W=0.445u L=180.00n
MM42 net0163 SE net0155 VPW n18 W=0.445u L=180.00n
MM47 SEN SE VSS VPW n18 W=0.52u L=180.00n
MM37 net100 cn net0264 VPW n18 W=0.42u L=180.00n
MM38 net0264 SDN net0260 VPW n18 W=0.42u L=180.00n
MM33 net108 c net0292 VPW n18 W=0.445u L=180.00n
MM45 net0163 cn net108 VPW n18 W=0.445u L=180.00n
MM31 net0276 net108 VSS VPW n18 W=0.49u L=180.00n
MM28 net0163 D net0320 VPW n18 W=0.445u L=180.00n
MM39 net0260 net112 VSS VPW n18 W=0.42u L=180.00n
MM1 net0320 SEN VSS VPW n18 W=0.445u L=180.00n
MM7 cn c VSS VPW n18 W=420.00n L=180.00n
MM3 c CKN VSS VPW n18 W=250.00n L=180.00n
MM19 net112 net100 net77 VPW n18 W=0.53u L=180.00n
MM18 net77 RDN VSS VPW n18 W=0.53u L=180.00n
MM23 net0292 RDN net93 VPW n18 W=0.445u L=180.00n
MM22 net93 net101 VSS VPW n18 W=0.445u L=180.00n
MM15 net101 c net100 VPW n18 W=0.42u L=180.00n
MM12 net101 SDN net0276 VPW n18 W=0.49u L=180.00n
MM4 Q net112 VSS VPW n18 W=0.72u L=180.00n
.ENDS SNDSRNQUHDV1
.SUBCKT SNDSRNQUHDV2 CKN D Q RDN SDN SE SI VDD VSS VNW VPW
MM40 net0163 SEN net082 VNW p18 W=0.36u L=180.00n
MM29 net0163 D net61 VNW p18 W=0.69u L=180.00n
MM41 net082 SI VDD VNW p18 W=0.36u L=180.00n
MM46 SEN SE VDD VNW p18 W=0.485u L=180.00n
MM44 net0163 c net108 VNW p18 W=0.42u L=180.00n
MM30 net101 SDN VDD VNW p18 W=0.37u L=180.00n
MM32 net108 cn net88 VNW p18 W=0.42u L=180.00n
MM21 net88 net101 VDD VNW p18 W=0.42u L=180.00n
MM20 net88 RDN VDD VNW p18 W=0.42u L=180.00n
MM14 net101 cn net100 VNW p18 W=0.425u L=180.00n
MM10 net101 net108 VDD VNW p18 W=0.42u L=180.00n
MM6 cn c VDD VNW p18 W=250.00n L=180.00n
MM2 c CKN VDD VNW p18 W=420.00n L=180.00n
MM0 net61 SE VDD VNW p18 W=0.69u L=180.00n
MM16 net112 RDN VDD VNW p18 W=0.42u L=180.00n
MM17 net112 net100 VDD VNW p18 W=0.42u L=180.00n
MM5 Q net112 VDD VNW p18 W=2.02u L=180.00n
MM34 net0204 net112 VDD VNW p18 W=0.42u L=180.00n
MM35 net0204 SDN VDD VNW p18 W=0.42u L=180.00n
MM36 net100 c net0204 VNW p18 W=0.425u L=180.00n
MM43 net0155 SI VSS VPW n18 W=0.445u L=180.00n
MM42 net0163 SE net0155 VPW n18 W=0.445u L=180.00n
MM47 SEN SE VSS VPW n18 W=0.52u L=180.00n
MM37 net100 cn net0264 VPW n18 W=0.42u L=180.00n
MM38 net0264 SDN net0260 VPW n18 W=0.42u L=180.00n
MM33 net108 c net0292 VPW n18 W=0.445u L=180.00n
MM45 net0163 cn net108 VPW n18 W=0.445u L=180.00n
MM31 net0276 net108 VSS VPW n18 W=0.49u L=180.00n
MM28 net0163 D net0320 VPW n18 W=0.445u L=180.00n
MM39 net0260 net112 VSS VPW n18 W=0.42u L=180.00n
MM1 net0320 SEN VSS VPW n18 W=0.445u L=180.00n
MM7 cn c VSS VPW n18 W=420.00n L=180.00n
MM3 c CKN VSS VPW n18 W=250.00n L=180.00n
MM19 net112 net100 net77 VPW n18 W=0.53u L=180.00n
MM18 net77 RDN VSS VPW n18 W=0.53u L=180.00n
MM23 net0292 RDN net93 VPW n18 W=0.445u L=180.00n
MM22 net93 net101 VSS VPW n18 W=0.445u L=180.00n
MM15 net101 c net100 VPW n18 W=0.42u L=180.00n
MM12 net101 SDN net0276 VPW n18 W=0.49u L=180.00n
MM4 Q net112 VSS VPW n18 W=1.4u L=180.00n
.ENDS SNDSRNQUHDV2
.SUBCKT TBUFUHDV0P7 I OE Z VDD VSS VNW VPW
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM3 net20 oen VSS VPW n18 W=430.00n L=180.00n
MM2 net20 OE net40 VPW n18 W=430.00n L=180.00n
MM4 Z net20 VSS VPW n18 W=560.00n L=180.00n
MM6 net20 I VSS VPW n18 W=430.00n L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM1 net20 oen net40 VNW p18 W=500.0n L=180.00n
MM0 net40 OE VDD VNW p18 W=400.0n L=180.00n
MM5 Z net40 VDD VNW p18 W=790.0n L=180.00n
MM7 net40 I VDD VNW p18 W=500.0n L=180.00n
.ENDS TBUFUHDV0P7
.SUBCKT TBUFUHDV1 I OE Z VDD VSS VNW VPW
MM7 net23 I VDD VNW p18 W=580.0n L=180.00n
MM0 net23 OE VDD VNW p18 W=400.0n L=180.00n
MM5 Z net23 VDD VNW p18 W=0.945u L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM1 net20 oen net23 VNW p18 W=500.0n L=180.00n
MM6 net20 I VSS VPW n18 W=430.00n L=180.00n
MM3 net20 oen VSS VPW n18 W=430.00n L=180.00n
MM4 Z net20 VSS VPW n18 W=0.56u L=180.00n
MM2 net20 OE net23 VPW n18 W=430.00n L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
.ENDS TBUFUHDV1
.SUBCKT TBUFUHDV12 I OE Z VDD VSS VNW VPW
MM1 net4 oen net7 VNW p18 W=0.79u L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM5 Z net7 VDD VNW p18 W=12.01u L=180.00n
MM0 net7 OE VDD VNW p18 W=790.0n L=180.00n
MM7 net7 I VDD VNW p18 W=4.04u L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM2 net4 OE net7 VPW n18 W=560.00n L=180.00n
MM4 Z net4 VSS VPW n18 W=7.92u L=180.00n
MM3 net4 oen VSS VPW n18 W=560.00n L=180.00n
MM6 net4 I VSS VPW n18 W=2.88u L=180.00n
.ENDS TBUFUHDV12
.SUBCKT TBUFUHDV16 I OE Z VDD VSS VNW VPW
MM6 net40 I VSS VPW n18 W=4.26u L=180.00n
MM3 net40 oen VSS VPW n18 W=630.00n L=180.00n
MM4 Z net40 VSS VPW n18 W=10.56u L=180.00n
MM2 net40 OE net43 VPW n18 W=560.00n L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM7 net43 I VDD VNW p18 W=5.99u L=180.00n
MM0 net43 OE VDD VNW p18 W=0.79u L=180.00n
MM5 Z net43 VDD VNW p18 W=16.02u L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM1 net40 oen net43 VNW p18 W=0.79u L=180.00n
.ENDS TBUFUHDV16
.SUBCKT TBUFUHDV2 I OE Z VDD VSS VNW VPW
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM2 net24 OE net27 VPW n18 W=430.00n L=180.00n
MM4 Z net24 VSS VPW n18 W=1.32u L=180.00n
MM3 net24 oen VSS VPW n18 W=430.00n L=180.00n
MM6 net24 I VSS VPW n18 W=630.00n L=180.00n
MM1 net24 oen net27 VNW p18 W=580.0n L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM5 Z net27 VDD VNW p18 W=1.96u L=180.00n
MM0 net27 OE VDD VNW p18 W=400.0n L=180.00n
MM7 net27 I VDD VNW p18 W=0.89u L=180.00n
.ENDS TBUFUHDV2
.SUBCKT TBUFUHDV24 I OE Z VDD VSS VNW VPW
MM6 net40 I VSS VPW n18 W=5.76u L=180.00n
MM3 net40 oen VSS VPW n18 W=720.00n L=180.00n
MM4 Z net40 VSS VPW n18 W=15.84u L=180.00n
MM2 net40 OE net43 VPW n18 W=1.39u L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM7 net43 I VDD VNW p18 W=8.08u L=180.00n
MM0 net43 OE VDD VNW p18 W=0.79u L=180.00n
MM5 Z net43 VDD VNW p18 W=24.03u L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM1 net40 oen net43 VNW p18 W=1.85u L=180.00n
.ENDS TBUFUHDV24
.SUBCKT TBUFUHDV3 I OE Z VDD VSS VNW VPW
MM6 net40 I VSS VPW n18 W=720.00n L=180.00n
MM3 net40 oen VSS VPW n18 W=430.00n L=180.00n
MM4 Z net40 VSS VPW n18 W=1.98u L=180.00n
MM2 net40 OE net43 VPW n18 W=430.00n L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM7 net43 I VDD VNW p18 W=1.01u L=180.00n
MM0 net43 OE VDD VNW p18 W=400.0n L=180.00n
MM5 Z net43 VDD VNW p18 W=2.97u L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM1 net40 oen net43 VNW p18 W=580.0n L=180.00n
.ENDS TBUFUHDV3
.SUBCKT TBUFUHDV4 I OE Z VDD VSS VNW VPW
MM1 net4 oen net7 VNW p18 W=580.0n L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM5 Z net7 VDD VNW p18 W=3.98u L=180.00n
MM0 net7 OE VDD VNW p18 W=400.0n L=180.00n
MM7 net7 I VDD VNW p18 W=1.49u L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM2 net4 OE net7 VPW n18 W=430.00n L=180.00n
MM4 Z net4 VSS VPW n18 W=2.64u L=180.00n
MM3 net4 oen VSS VPW n18 W=430.00n L=180.00n
MM6 net4 I VSS VPW n18 W=1060.00n L=180.00n
.ENDS TBUFUHDV4
.SUBCKT TBUFUHDV6 I OE Z VDD VSS VNW VPW
MM6 net40 I VSS VPW n18 W=1.44u L=180.00n
MM3 net40 oen VSS VPW n18 W=430.00n L=180.00n
MM4 Z net40 VSS VPW n18 W=3.96u L=180.00n
MM2 net40 OE net43 VPW n18 W=430.00n L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM7 net43 I VDD VNW p18 W=2.02u L=180.00n
MM0 net43 OE VDD VNW p18 W=0.42u L=180.00n
MM5 Z net43 VDD VNW p18 W=6u L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM1 net40 oen net43 VNW p18 W=0.61u L=180.00n
.ENDS TBUFUHDV6
.SUBCKT TBUFUHDV8 I OE Z VDD VSS VNW VPW
MM1 net4 oen net7 VNW p18 W=790.00n L=180.00n
MM9 oen OE VDD VNW p18 W=0.49u L=180.00n
MM5 Z net7 VDD VNW p18 W=8.01u L=180.00n
MM0 net7 OE VDD VNW p18 W=500.0n L=180.00n
MM7 net7 I VDD VNW p18 W=2.99u L=180.00n
MM8 oen OE VSS VPW n18 W=430.00n L=180.00n
MM2 net4 OE net7 VPW n18 W=560.00n L=180.00n
MM4 Z net4 VSS VPW n18 W=5.28u L=180.00n
MM3 net4 oen VSS VPW n18 W=0.56u L=180.00n
MM6 net4 I VSS VPW n18 W=2.13u L=180.00n
.ENDS TBUFUHDV8
.SUBCKT XNOR2UHDV0P4 A1 A2 ZN VDD VSS VNW VPW
MM7 ZN A1 net8 VPW n18 W=0.28u L=180.00n
MM4 net8 a2n VSS VPW n18 W=0.28u L=180.00n
MM13 a2n a1n ZN VPW n18 W=0.28u L=180.00n
MM3 a1n A1 VSS VPW n18 W=0.28u L=180.00n
MM0 a2n A2 VSS VPW n18 W=0.28u L=180.00n
MM6 ZN a1n net27 VNW p18 W=490.0n L=180.00n
MM5 net27 a2n VDD VNW p18 W=490.0n L=180.00n
MM11 a2n A1 ZN VNW p18 W=490.0n L=180.00n
MM2 a1n A1 VDD VNW p18 W=490.0n L=180.00n
MM1 a2n A2 VDD VNW p18 W=490.0n L=180.00n
.ENDS XNOR2UHDV0P4
.SUBCKT XNOR2UHDV0P7 A1 A2 ZN VDD VSS VNW VPW
MM5 net60 a2n VDD VNW p18 W=790.0n L=180.00n
MM6 ZN a1n net60 VNW p18 W=790.0n L=180.00n
MM2 a1n A1 VDD VNW p18 W=790.0n L=180.00n
MM11 a2n A1 ZN VNW p18 W=790.0n L=180.00n
MM1 a2n A2 VDD VNW p18 W=790.0n L=180.00n
MM7 ZN A1 net73 VPW n18 W=540.00n L=180.00n
MM4 net73 a2n VSS VPW n18 W=540.00n L=180.00n
MM13 a2n a1n ZN VPW n18 W=540.00n L=180.00n
MM3 a1n A1 VSS VPW n18 W=540.00n L=180.00n
MM0 a2n A2 VSS VPW n18 W=540.00n L=180.00n
.ENDS XNOR2UHDV0P7
.SUBCKT XNOR2UHDV1 A1 A2 ZN VDD VSS VNW VPW
MM6 ZN a1n net60 VNW p18 W=0.925u L=180.00n
MM5 net60 a2n VDD VNW p18 W=0.925u L=180.00n
MM11 a2n A1 ZN VNW p18 W=0.95u L=180.00n
MM2 a1n A1 VDD VNW p18 W=0.95u L=180.00n
MM1 a2n A2 VDD VNW p18 W=0.58u L=180.00n
MM0 a2n A2 VSS VPW n18 W=720.00n L=180.00n
MM3 a1n A1 VSS VPW n18 W=720.00n L=180.00n
MM7 ZN A1 net73 VPW n18 W=720.00n L=180.00n
MM4 net73 a2n VSS VPW n18 W=720.00n L=180.00n
MM13 a2n a1n ZN VPW n18 W=720.00n L=180.00n
.ENDS XNOR2UHDV1
.SUBCKT XNOR2UHDV2 A1 A2 ZN VDD VSS VNW VPW
MM6 net65 a2n VDD VNW p18 W=0.925u L=180.00n
MM11 net65 a1n ZN VNW p18 W=0.925u L=180.00n
MM2 a1n A1 VDD VNW p18 W=2.02u L=180.00n
MM1 a2n A2 VDD VNW p18 W=2.02u L=180.00n
MM4 a2n A1 ZN VNW p18 W=0.925u L=180.00n
MM7 net65 a2n VSS VPW n18 W=0.72u L=180.00n
MM3 a1n A1 VSS VPW n18 W=1.44u L=180.00n
MM13 net65 A1 ZN VPW n18 W=690.00n L=180.00n
MM0 a2n A2 VSS VPW n18 W=1.44u L=180.00n
MM5 a2n a1n ZN VPW n18 W=740.00n L=180.00n
.ENDS XNOR2UHDV2
.SUBCKT XNOR2UHDV4 A1 A2 ZN VDD VSS VNW VPW
MM7 net57 a2n VSS VPW n18 W=720.00n L=180.00n
MM3 a1n A1 VSS VPW n18 W=2.88u L=180.00n
MM13 net57 A1 ZN VPW n18 W=2.24u L=180.00n
MM0 a2n A2 VSS VPW n18 W=2.88u L=180.00n
MM5 a2n a1n ZN VPW n18 W=2.33u L=180.00n
MM11 net57 a1n ZN VNW p18 W=2.775u L=180.00n
MM2 a1n A1 VDD VNW p18 W=4.04u L=180.00n
MM1 a2n A2 VDD VNW p18 W=4.04u L=180.00n
MM4 a2n A1 ZN VNW p18 W=3.35u L=180.00n
MM6 net57 a2n VDD VNW p18 W=1.01u L=180.00n
.ENDS XNOR2UHDV4
.SUBCKT XNOR3UHDV0P7 A1 A2 A3 ZN VDD VSS VNW VPW
MM14 ZN net56 VDD VNW p18 W=790.0n L=180.00n
MM18 net49 net81 VDD VNW p18 W=500.0n L=180.00n
MM8 net61 A3 net56 VNW p18 W=500.0n L=180.00n
MM7 net72 a3n net56 VNW p18 W=0.495u L=180.00n
MM17 net61 net72 VDD VNW p18 W=500.0n L=180.00n
MM11 net81 A2 net72 VNW p18 W=500.0n L=180.00n
MM10 net49 a2n net72 VNW p18 W=500.0n L=180.00n
MM2 a2n A2 VDD VNW p18 W=500.0n L=180.00n
MM4 a3n A3 VDD VNW p18 W=500.0n L=180.00n
MM1 net81 A1 VDD VNW p18 W=500.0n L=180.00n
MM15 ZN net56 VSS VPW n18 W=560.00n L=180.00n
MM19 net49 net81 VSS VPW n18 W=430.00n L=180.00n
MM9 net61 a3n net56 VPW n18 W=430.00n L=180.00n
MM6 net72 A3 net56 VPW n18 W=430.00n L=180.00n
MM16 net61 net72 VSS VPW n18 W=430.00n L=180.00n
MM13 net81 a2n net72 VPW n18 W=360.00n L=180.00n
MM12 net49 A2 net72 VPW n18 W=430.00n L=180.00n
MM3 a2n A2 VSS VPW n18 W=430.00n L=180.00n
MM5 a3n A3 VSS VPW n18 W=430.00n L=180.00n
MM0 net81 A1 VSS VPW n18 W=360.00n L=180.00n
.ENDS XNOR3UHDV0P7
.SUBCKT XNOR3UHDV1 A1 A2 A3 ZN VDD VSS VNW VPW
MM16 net142 net109 VSS VPW n18 W=430.00n L=180.00n
MM15 ZN net137 VSS VPW n18 W=720.00n L=180.00n
MM9 net142 a3n net137 VPW n18 W=430.00n L=180.00n
MM6 net109 A3 net137 VPW n18 W=430.00n L=180.00n
MM0 net126 A1 VSS VPW n18 W=360.00n L=180.00n
MM3 a2n A2 VSS VPW n18 W=430.00n L=180.00n
MM5 a3n A3 VSS VPW n18 W=430.00n L=180.00n
MM19 net114 net126 VSS VPW n18 W=430.00n L=180.00n
MM13 net126 a2n net109 VPW n18 W=360.00n L=180.00n
MM12 net114 A2 net109 VPW n18 W=430.00n L=180.00n
MM17 net142 net109 VDD VNW p18 W=580.0n L=180.00n
MM14 ZN net137 VDD VNW p18 W=1.01u L=180.00n
MM8 net142 A3 net137 VNW p18 W=580.0n L=180.00n
MM7 net109 a3n net137 VNW p18 W=0.495u L=180.00n
MM1 net126 A1 VDD VNW p18 W=580.0n L=180.00n
MM2 a2n A2 VDD VNW p18 W=580.0n L=180.00n
MM4 a3n A3 VDD VNW p18 W=0.57u L=180.00n
MM18 net114 net126 VDD VNW p18 W=580.0n L=180.00n
MM11 net126 A2 net109 VNW p18 W=580.0n L=180.00n
MM10 net114 a2n net109 VNW p18 W=580.0n L=180.00n
.ENDS XNOR3UHDV1
.SUBCKT XNOR3UHDV2 A1 A2 A3 ZN VDD VSS VNW VPW
MM16 net142 net109 VSS VPW n18 W=0.675u L=180.00n
MM15 ZN net137 VSS VPW n18 W=1.44u L=180.00n
MM9 net142 a3n net137 VPW n18 W=0.675u L=180.00n
MM6 net109 A3 net137 VPW n18 W=0.615u L=180.00n
MM0 net126 A1 VSS VPW n18 W=690.00n L=180.00n
MM3 a2n A2 VSS VPW n18 W=0.675u L=180.00n
MM5 a3n A3 VSS VPW n18 W=0.66u L=180.00n
MM19 net114 net126 VSS VPW n18 W=690.00n L=180.00n
MM13 net126 a2n net109 VPW n18 W=690.00n L=180.00n
MM12 net114 A2 net109 VPW n18 W=690.00n L=180.00n
MM17 net142 net109 VDD VNW p18 W=950.0n L=180.00n
MM14 ZN net137 VDD VNW p18 W=2.02u L=180.00n
MM8 net142 A3 net137 VNW p18 W=0.925u L=180.00n
MM7 net109 a3n net137 VNW p18 W=0.925u L=180.00n
MM1 net126 A1 VDD VNW p18 W=950.0n L=180.00n
MM2 a2n A2 VDD VNW p18 W=0.865u L=180.00n
MM4 a3n A3 VDD VNW p18 W=0.925u L=180.00n
MM18 net114 net126 VDD VNW p18 W=950.0n L=180.00n
MM11 net126 A2 net109 VNW p18 W=0.865u L=180.00n
MM10 net114 a2n net109 VNW p18 W=0.925u L=180.00n
.ENDS XNOR3UHDV2
.SUBCKT XOR2UHDV0P4 A1 A2 Z VDD VSS VNW VPW
MM1 a2n A2 VDD VNW p18 W=490.0n L=180.00n
MM2 a1n A1 VDD VNW p18 W=490.0n L=180.00n
MM11 a2n a1n Z VNW p18 W=490.0n L=180.00n
MM5 net23 a2n VDD VNW p18 W=490.0n L=180.00n
MM6 Z A1 net23 VNW p18 W=490.0n L=180.00n
MM0 a2n A2 VSS VPW n18 W=0.28u L=180.00n
MM3 a1n A1 VSS VPW n18 W=0.28u L=180.00n
MM13 a2n A1 Z VPW n18 W=0.28u L=180.00n
MM4 net36 a2n VSS VPW n18 W=0.28u L=180.00n
MM7 Z a1n net36 VPW n18 W=0.28u L=180.00n
.ENDS XOR2UHDV0P4
.SUBCKT XOR2UHDV0P7 A1 A2 Z VDD VSS VNW VPW
MM0 a2n A2 VSS VPW n18 W=560.00n L=180.00n
MM3 a1n A1 VSS VPW n18 W=560.00n L=180.00n
MM13 a2n A1 Z VPW n18 W=560.00n L=180.00n
MM4 net45 a2n VSS VPW n18 W=560.00n L=180.00n
MM7 Z a1n net45 VPW n18 W=560.00n L=180.00n
MM1 a2n A2 VDD VNW p18 W=790.0n L=180.00n
MM2 a1n A1 VDD VNW p18 W=790.0n L=180.00n
MM11 a2n a1n Z VNW p18 W=790.0n L=180.00n
MM5 net64 a2n VDD VNW p18 W=790.0n L=180.00n
MM6 Z A1 net64 VNW p18 W=790.0n L=180.00n
.ENDS XOR2UHDV0P7
.SUBCKT XOR2UHDV1 A1 A2 Z VDD VSS VNW VPW
MM3 a1n A1 VSS VPW n18 W=720.00n L=180.00n
MM13 a2n A1 Z VPW n18 W=800.00n L=180.00n
MM4 net45 a2n VSS VPW n18 W=720.00n L=180.00n
MM7 Z a1n net45 VPW n18 W=0.72u L=180.00n
MM0 a2n A2 VSS VPW n18 W=720.00n L=180.00n
MM1 a2n A2 VDD VNW p18 W=1.01u L=180.00n
MM2 a1n A1 VDD VNW p18 W=1.01u L=180.00n
MM11 a2n a1n Z VNW p18 W=1170.0n L=180.00n
MM5 net64 a2n VDD VNW p18 W=1.01u L=180.00n
MM6 Z A1 net64 VNW p18 W=1.01u L=180.00n
.ENDS XOR2UHDV1
.SUBCKT XOR2UHDV2 A1 A2 Z VDD VSS VNW VPW
MM10 net77 a2n VDD VNW p18 W=0.925u L=180.00n
MM7 net77 A1 Z VNW p18 W=0.925u L=180.00n
MM11 a2n a1n Z VNW p18 W=0.925u L=180.00n
MM2 a1n A1 VDD VNW p18 W=2.02u L=180.00n
MM1 a2n A2 VDD VNW p18 W=2.02u L=180.00n
MM9 net77 a2n VSS VPW n18 W=0.72u L=180.00n
MM8 net77 a1n Z VPW n18 W=720.00n L=180.00n
MM13 a2n A1 Z VPW n18 W=720.00n L=180.00n
MM3 a1n A1 VSS VPW n18 W=1.37u L=180.00n
MM0 a2n A2 VSS VPW n18 W=1.44u L=180.00n
.ENDS XOR2UHDV2
.SUBCKT XOR2UHDV4 A1 A2 Z VDD VSS VNW VPW
MM1 a2n A2 VDD VNW p18 W=4.04u L=180.00n
MM2 a1n A1 VDD VNW p18 W=4.04u L=180.00n
MM11 a2n a1n Z VNW p18 W=3.33u L=180.00n
MM7 net40 A1 Z VNW p18 W=2.715u L=180.00n
MM10 net40 a2n VDD VNW p18 W=1.01u L=180.00n
MM0 a2n A2 VSS VPW n18 W=2.88u L=180.00n
MM3 a1n A1 VSS VPW n18 W=2.88u L=180.00n
MM13 a2n A1 Z VPW n18 W=2.33u L=180.00n
MM8 net40 a1n Z VPW n18 W=2.23u L=180.00n
MM9 net40 a2n VSS VPW n18 W=720.00n L=180.00n
.ENDS XOR2UHDV4
.SUBCKT XOR3UHDV0P7T A1 A2 A3 Z VDD VSS VNW VPW
MM0 net5 A1 VSS VPW n18 W=360.00n L=180.00n
MM5 a3n A3 VSS VPW n18 W=430.00n L=180.00n
MM3 a2n A2 VSS VPW n18 W=430.00n L=180.00n
MM12 net37 A2 net20 VPW n18 W=430.00n L=180.00n
MM13 net5 a2n net20 VPW n18 W=360.00n L=180.00n
MM16 net25 net20 VSS VPW n18 W=430.00n L=180.00n
MM6 net20 a3n net36 VPW n18 W=0.42u L=180.00n
MM9 net25 A3 net36 VPW n18 W=430.00n L=180.00n
MM19 net37 net5 VSS VPW n18 W=430.00n L=180.00n
MM15 Z net36 VSS VPW n18 W=560.00n L=180.00n
MM1 net5 A1 VDD VNW p18 W=500.0n L=180.00n
MM4 a3n A3 VDD VNW p18 W=500.0n L=180.00n
MM2 a2n A2 VDD VNW p18 W=500.0n L=180.00n
MM10 net37 a2n net20 VNW p18 W=500.0n L=180.00n
MM11 net5 A2 net20 VNW p18 W=500.0n L=180.00n
MM17 net25 net20 VDD VNW p18 W=500.0n L=180.00n
MM7 net20 A3 net36 VNW p18 W=500.0n L=180.00n
MM8 net25 a3n net36 VNW p18 W=500.0n L=180.00n
MM18 net37 net5 VDD VNW p18 W=500.0n L=180.00n
MM14 Z net36 VDD VNW p18 W=790.0n L=180.00n
.ENDS XOR3UHDV0P7T
.SUBCKT XOR3UHDV1T A1 A2 A3 Z VDD VSS VNW VPW
MM0 net5 A1 VSS VPW n18 W=360.00n L=180.00n
MM5 a3n A3 VSS VPW n18 W=430.00n L=180.00n
MM3 a2n A2 VSS VPW n18 W=430.00n L=180.00n
MM12 net37 A2 net20 VPW n18 W=430.00n L=180.00n
MM13 net5 a2n net20 VPW n18 W=360.00n L=180.00n
MM16 net25 net20 VSS VPW n18 W=430.00n L=180.00n
MM6 net20 a3n net36 VPW n18 W=340.00n L=180.00n
MM9 net25 A3 net36 VPW n18 W=430.00n L=180.00n
MM19 net37 net5 VSS VPW n18 W=430.00n L=180.00n
MM15 Z net36 VSS VPW n18 W=720.00n L=180.00n
MM1 net5 A1 VDD VNW p18 W=580.0n L=180.00n
MM4 a3n A3 VDD VNW p18 W=580.0n L=180.00n
MM2 a2n A2 VDD VNW p18 W=580.0n L=180.00n
MM10 net37 a2n net20 VNW p18 W=580.0n L=180.00n
MM11 net5 A2 net20 VNW p18 W=580.0n L=180.00n
MM17 net25 net20 VDD VNW p18 W=580.0n L=180.00n
MM7 net20 A3 net36 VNW p18 W=580.0n L=180.00n
MM8 net25 a3n net36 VNW p18 W=580.0n L=180.00n
MM18 net37 net5 VDD VNW p18 W=580.0n L=180.00n
MM14 Z net36 VDD VNW p18 W=990.0n L=180.00n
.ENDS XOR3UHDV1T
.SUBCKT XOR3UHDV2T A1 A2 A3 Z VDD VSS VNW VPW
MM18 net49 net81 VDD VNW p18 W=950.0n L=180.00n
MM17 net61 net72 VDD VNW p18 W=950.0n L=180.00n
MM14 Z net56 VDD VNW p18 W=2.02u L=180.00n
MM11 net81 A2 net72 VNW p18 W=0.865u L=180.00n
MM10 net49 a2n net72 VNW p18 W=0.925u L=180.00n
MM8 net61 a3n net56 VNW p18 W=0.925u L=180.00n
MM7 net72 A3 net56 VNW p18 W=0.865u L=180.00n
MM2 a2n A2 VDD VNW p18 W=0.865u L=180.00n
MM1 net81 A1 VDD VNW p18 W=950.0n L=180.00n
MM4 a3n A3 VDD VNW p18 W=0.865u L=180.00n
MM19 net49 net81 VSS VPW n18 W=690.00n L=180.00n
MM16 net61 net72 VSS VPW n18 W=0.675u L=180.00n
MM15 Z net56 VSS VPW n18 W=1.44u L=180.00n
MM13 net81 a2n net72 VPW n18 W=690.00n L=180.00n
MM12 net49 A2 net72 VPW n18 W=690.00n L=180.00n
MM9 net61 A3 net56 VPW n18 W=0.675u L=180.00n
MM3 a2n A2 VSS VPW n18 W=0.675u L=180.00n
MM0 net81 A1 VSS VPW n18 W=690.00n L=180.00n
MM6 net72 a3n net56 VPW n18 W=0.615u L=180.00n
MM5 a3n A3 VSS VPW n18 W=690.00n L=180.00n
.ENDS XOR3UHDV2T
